module ps7_axi_wrapper
(
  `ifdef USE_CAN0
    output wire CAN0_PHY_TX,
    input wire CAN0_PHY_RX,
  `endif

  `ifdef USE_CAN1
    output wire CAN1_PHY_TX,  
    input wire CAN1_PHY_RX,
  `endif

  // Ethernet wires
  `ifdef USE_ENET0
    output wire ENET0_GMII_TX_EN,
    output wire ENET0_GMII_TX_ER,
    output wire ENET0_MDIO_MDC,
    output wire ENET0_MDIO_O,
    output wire ENET0_MDIO_T,
    output wire ENET0_PTP_DELAY_REQ_RX,
    output wire ENET0_PTP_DELAY_REQ_TX,
    output wire ENET0_PTP_PDELAY_REQ_RX,
    output wire ENET0_PTP_PDELAY_REQ_TX,
    output wire ENET0_PTP_PDELAY_RESP_RX,
    output wire ENET0_PTP_PDELAY_RESP_TX,
    output wire ENET0_PTP_SYNC_FRAME_RX,
    output wire ENET0_PTP_SYNC_FRAME_TX,
    output wire ENET0_SOF_RX,
    output wire ENET0_SOF_TX,
    output wire [7:0] ENET0_GMII_TXD,  
    input wire ENET0_GMII_COL,
    input wire ENET0_GMII_CRS,
    input wire ENET0_GMII_RX_CLK,
    input wire ENET0_GMII_RX_DV,
    input wire ENET0_GMII_RX_ER,
    input wire ENET0_GMII_TX_CLK,
    input wire ENET0_MDIO_I,
    input wire ENET0_EXT_INTIN,
    input wire [7:0] ENET0_GMII_RXD,  
  `endif
  `ifdef USE_ENET1
    output wire ENET1_GMII_TX_EN,
    output wire ENET1_GMII_TX_ER,
    output wire ENET1_MDIO_MDC,
    output wire ENET1_MDIO_O,
    output wire ENET1_MDIO_T,
    output wire ENET1_PTP_DELAY_REQ_RX,
    output wire ENET1_PTP_DELAY_REQ_TX,
    output wire ENET1_PTP_PDELAY_REQ_RX,
    output wire ENET1_PTP_PDELAY_REQ_TX,
    output wire ENET1_PTP_PDELAY_RESP_RX,
    output wire ENET1_PTP_PDELAY_RESP_TX,
    output wire ENET1_PTP_SYNC_FRAME_RX,
    output wire ENET1_PTP_SYNC_FRAME_TX,
    output wire ENET1_SOF_RX,
    output wire ENET1_SOF_TX,
    output wire [7:0] ENET1_GMII_TXD,  
    input wire ENET1_GMII_COL,
    input wire ENET1_GMII_CRS,
    input wire ENET1_GMII_RX_CLK,
    input wire ENET1_GMII_RX_DV,
    input wire ENET1_GMII_RX_ER,
    input wire ENET1_GMII_TX_CLK,
    input wire ENET1_MDIO_I,
    input wire ENET1_EXT_INTIN,
    input wire [7:0] ENET1_GMII_RXD,  
  `endif

  // 4 DMA ports
  `ifdef USE_DMA0
    input wire DMA0_ACLK,
    output wire DMA0_RESET,
    output wire [1:0] DMA0_DATYPE,  
    input wire [1:0] DMA0_DRTYPE,
    output wire DMA0_DAVALID,
    output wire DMA0_DRREADY,
    input wire DMA0_DAREADY,
    input wire DMA0_DRLAST,
    input wire DMA0_DRVALID,
  `endif
  `ifdef USE_DMA1
    input wire DMA1_ACLK,
    output wire DMA1_RESET,
    output wire [1:0] DMA1_DATYPE,  
    input wire [1:0] DMA1_DRTYPE,
    output wire DMA1_DAVALID,
    output wire DMA1_DRREADY,
    input wire DMA1_DAREADY,
    input wire DMA1_DRLAST,
    input wire DMA1_DRVALID,
  `endif
  `ifdef USE_DMA2
    input wire DMA2_ACLK,
    output wire DMA2_RESET,  
    output wire [1:0] DMA2_DATYPE,  
    input wire [1:0] DMA2_DRTYPE,
    output wire DMA2_DAVALID,
    output wire DMA2_DRREADY,
    input wire DMA2_DAREADY,
    input wire DMA2_DRLAST,
    input wire DMA2_DRVALID,
  `endif
  `ifdef USE_DMA3
    input wire DMA3_ACLK,
    output wire DMA3_RESET,  
    output wire [1:0] DMA3_DATYPE,    
    input wire [1:0] DMA3_DRTYPE,
    output wire DMA3_DRREADY,
    input wire DMA3_DAREADY,
    input wire DMA3_DRLAST,
    input wire DMA3_DRVALID,  
    output wire DMA3_DAVALID,
  `endif

  // tristate GPIO wires + 54 MIO
  `ifdef USE_GPIO
    input wire [63:0] GPIO_I,
    output wire [63:0] GPIO_O,
    output wire [63:0] GPIO_T,
  `endif
  `ifdef USE_MIO
    inout wire [53:0] MIO,
  `endif

  // 2x I2C buses
  `ifdef USE_I2C0
    input wire I2C0_SDA_I,
    output wire I2C0_SDA_O,
    output wire I2C0_SDA_T,
    input wire I2C0_SCL_I,
    output wire I2C0_SCL_O,
    output wire I2C0_SCL_T,
  `endif
  `ifdef USE_I2C1
    input wire I2C1_SDA_I,
    output wire I2C1_SDA_O,
    output wire I2C1_SDA_T,
    input wire I2C1_SCL_I,
    output wire I2C1_SCL_O,
    output wire I2C1_SCL_T,
  `endif

  // 2x SDIO 
  `ifdef USE_SDIO0
    output wire SDIO0_CLK,
    input wire SDIO0_CLK_FB,
    output wire SDIO0_CMD_O,
    input wire SDIO0_CMD_I,
    output wire SDIO0_CMD_T,
    input wire [3:0] SDIO0_DATA_I,
    output wire [3:0] SDIO0_DATA_O,
    output wire [3:0] SDIO0_DATA_T,
    output wire SDIO0_LED,
    input wire SDIO0_CDN,
    input wire SDIO0_WP,  
    output wire SDIO0_BUSPOW,
    output wire [2:0] SDIO0_BUSVOLT,
  `endif
  `ifdef USE_SDIO1
    output wire SDIO1_CLK,
    input wire SDIO1_CLK_FB,
    output wire SDIO1_CMD_O,
    input wire SDIO1_CMD_I,
    output wire SDIO1_CMD_T,
    input wire [3:0] SDIO1_DATA_I,
    output wire [3:0] SDIO1_DATA_O,
    output wire [3:0] SDIO1_DATA_T,
    output wire SDIO1_LED,
    input wire SDIO1_CDN,
    input wire SDIO1_WP,
    output wire SDIO1_BUSPOW,
    output wire [2:0] SDIO1_BUSVOLT,
  `endif

  // 2x SPI
  `ifdef USE_SPI0
    input wire SPI0_SCLK_I,
    output  wire SPI0_SCLK_O,
    output wire SPI0_SCLK_T,
    input wire SPI0_MOSI_I,
    output wire SPI0_MOSI_O,
    output wire SPI0_MOSI_T,
    input wire SPI0_MISO_I,
    output wire SPI0_MISO_O,
    output wire SPI0_MISO_T,
    input wire SPI0_SS_I,
    output wire SPI0_SS_O,
    output wire SPI0_SS1_O,
    output wire SPI0_SS2_O,
    output wire SPI0_SS_T,
  `endif
  `ifdef USE_SPI1
    input wire SPI1_SCLK_I,
    output wire SPI1_SCLK_O,
    output wire SPI1_SCLK_T,
    input wire SPI1_MOSI_I,
    output wire SPI1_MOSI_O,
    output wire SPI1_MOSI_T,
    input wire SPI1_MISO_I,
    output wire SPI1_MISO_O,
    output wire SPI1_MISO_T,
    input wire SPI1_SS_I,
    output wire SPI1_SS_O,
    output wire SPI1_SS1_O,
    output wire SPI1_SS2_O,
    output wire SPI1_SS_T,
  `endif
  // 2 x UART
  `ifdef USE_UART0
    output wire UART0_DTRN,
    output wire UART0_RTSN, 
    output wire UART0_TX,
    input wire UART0_CTSN,
    input wire UART0_DCDN,
    input wire UART0_DSRN,
    input wire UART0_RIN,
    input wire UART0_RX,
  `endif
  `ifdef USE_UART1
    output wire UART1_DTRN,
    output wire UART1_RTSN,  
    output wire UART1_TX,
    input wire UART1_CTSN,
    input wire UART1_DCDN,
    input wire UART1_DSRN,
    input wire UART1_RIN,
    input wire UART1_RX,
  `endif

  // trace, debug and jtag
  `ifdef USE_JTAG
    input wire PJTAG_TCK,
    input wire PJTAG_TMS,
    input wire PJTAG_TDI,
    output wire PJTAG_TDO,
  `endif
  `ifdef USE_TTC0
    output wire TTC0_WAVE0_OUT,
    output wire TTC0_WAVE1_OUT,
    output wire TTC0_WAVE2_OUT,
    input wire TTC0_CLK0_IN,
    input wire TTC0_CLK1_IN,
    input wire TTC0_CLK2_IN,
  `endif
  `ifdef USE_TTC1
  output wire TTC1_WAVE0_OUT,
  output wire TTC1_WAVE1_OUT,
  output wire TTC1_WAVE2_OUT,
  input wire TTC1_CLK0_IN,
  input wire TTC1_CLK1_IN,
  input wire TTC1_CLK2_IN,
  `endif
  `ifdef USE_TRACE
    input wire TRACE_CLK,
    output wire TRACE_CTL,
    output wire [31:0] TRACE_DATA,
    output wire TRACE_CLK_OUT,

    input wire [31:0] FTMD_TRACEIN_DATA,
    input wire FTMD_TRACEIN_VALID,
    input wire FTMD_TRACEIN_CLK,
    input wire [3:0]  FTMD_TRACEIN_ATID,
    input wire FTMT_F2P_TRIG_0,
    output wire FTMT_F2P_TRIGACK_0,
    input wire FTMT_F2P_TRIG_1,
    output wire FTMT_F2P_TRIGACK_1,
    input wire FTMT_F2P_TRIG_2,
    output wire FTMT_F2P_TRIGACK_2,
    input wire FTMT_F2P_TRIG_3,
    output wire FTMT_F2P_TRIGACK_3,
    input wire [31:0] FTMT_F2P_DEBUG,
    input wire FTMT_P2F_TRIGACK_0,
    output wire FTMT_P2F_TRIG_0,
    input wire FTMT_P2F_TRIGACK_1,
    output wire FTMT_P2F_TRIG_1,
    input wire FTMT_P2F_TRIGACK_2,
    output wire FTMT_P2F_TRIG_2,
    input wire FTMT_P2F_TRIGACK_3,
    output wire FTMT_P2F_TRIG_3,
    output wire [31:0] FTMT_P2F_DEBUG,
  `endif
  `ifdef USE_WATCHDOG
    input wire WDT_CLK_IN,
    output wire WDT_RST_OUT,
  `endif
  `ifdef USE_USB0
    output wire [1:0] USB0_PORT_INDCTL,
    output wire USB0_VBUS_PWRSELECT,
    input wire USB0_VBUS_PWRFAULT,
  `endif
  `ifdef USE_USB1
    output wire [1:0]  USB1_PORT_INDCTL,
    output wire USB1_VBUS_PWRSELECT,
    input wire USB1_VBUS_PWRFAULT,
  `endif

  `ifdef USE_INTERRUPTS
    // events and interrupts
    output wire IRQ_P2F_DMAC_ABORT,
    output wire IRQ_P2F_DMAC0,
    output wire IRQ_P2F_DMAC1,
    output wire IRQ_P2F_DMAC2,
    output wire IRQ_P2F_DMAC3,
    output wire IRQ_P2F_DMAC4,
    output wire IRQ_P2F_DMAC5,
    output wire IRQ_P2F_DMAC6,
    output wire IRQ_P2F_DMAC7,
    output wire IRQ_P2F_SMC,
    output wire IRQ_P2F_QSPI,
    output wire IRQ_P2F_CTI,
    output wire IRQ_P2F_GPIO,
    output wire IRQ_P2F_USB0,
    output wire IRQ_P2F_ENET0,
    output wire IRQ_P2F_ENET_WAKE0,
    output wire IRQ_P2F_SDIO0,
    output wire IRQ_P2F_I2C0,
    output wire IRQ_P2F_SPI0,
    output wire IRQ_P2F_UART0,
    output wire IRQ_P2F_CAN0,
    output wire IRQ_P2F_USB1,
    output wire IRQ_P2F_ENET1,
    output wire IRQ_P2F_ENET_WAKE1,
    output wire IRQ_P2F_SDIO1,
    output wire IRQ_P2F_I2C1,
    output wire IRQ_P2F_SPI1,
    output wire IRQ_P2F_UART1,
    output wire IRQ_P2F_CAN1,
    input  wire Core0_nFIQ,
    input  wire Core0_nIRQ,
    input  wire Core1_nFIQ,
    input  wire Core1_nIRQ,
    input  wire [15:0] IRQ_F2P,
    input wire SRAM_INTIN,
  `endif
  `ifdef USE_PS_EVENTS
    output wire EVENT_EVENTO,
    input wire EVENT_EVENTI,   
    output wire [1:0] EVENT_STANDBYWFE,
    output wire [1:0] EVENT_STANDBYWFI,
  `endif
  `ifdef USE_FPGA_IDLE
    input wire FPGA_IDLE,
  `endif

  // 4 frabric clks
  `ifdef USE_FCLK0
    output wire FCLK0_CLK,
    output wire FCLK0_RESET,
  `endif
  `ifdef USE_FCLK1
    output wire FCLK1_CLK,
    output wire FCLK1_RESET,
  `endif
  `ifdef USE_FCLK2
    output wire FCLK2_CLK,
    output wire FCLK2_RESET,
  `endif
  `ifdef USE_FCLK3
    output wire FCLK3_CLK,
    output wire FCLK3_RESET,
  `endif

  // AXI3+ (3 with some optional Axi4 wires)
  // direction is from PS point of view
  // 2 PS Master General Purpose ports
  // 2 PS Slave General Purpose ports
  // 1 PS Slave ACP port
  // 4 PS Slave High Performance ports

  `ifdef PS_MASTER_AXI_GP0
    //M_AXI_GP0  
    input wire M_AXI_GP0_clk,
    output wire M_AXI_GP0_reset,

    output wire M_AXI_GP0_ar_valid,
    output wire M_AXI_GP0_aw_valid,
    input wire M_AXI_GP0_r_valid,
    output wire M_AXI_GP0_w_valid,
    input wire M_AXI_GP0_b_valid,

    input wire M_AXI_GP0_ar_ready,
    input wire M_AXI_GP0_aw_ready,
    output wire M_AXI_GP0_r_ready,
    input wire M_AXI_GP0_w_ready,
    output wire M_AXI_GP0_b_ready,

    output wire [31:0] M_AXI_GP0_ar_payload_addr,
    output wire [11:0] M_AXI_GP0_ar_payload_id,
    output wire [1:0] M_AXI_GP0_ar_payload_burst,
    output wire M_AXI_GP0_ar_payload_lock,
    output wire [2:0] M_AXI_GP0_ar_payload_size,
    output wire [2:0] M_AXI_GP0_ar_payload_prot,
    output wire [3:0] M_AXI_GP0_ar_payload_cache,
    output wire [7:0] M_AXI_GP0_ar_payload_len,
    output wire [3:0] M_AXI_GP0_ar_payload_qos,
    output wire [31:0] M_AXI_GP0_aw_payload_addr,
    output wire [11:0] M_AXI_GP0_aw_payload_id,
    output wire [1:0] M_AXI_GP0_aw_payload_burst,
    output wire M_AXI_GP0_aw_payload_lock,
    output wire [2:0] M_AXI_GP0_aw_payload_size,
    output wire [2:0] M_AXI_GP0_aw_payload_prot,
    output wire [3:0] M_AXI_GP0_aw_payload_cache,
    output wire [7:0] M_AXI_GP0_aw_payload_len,
    output wire [3:0] M_AXI_GP0_aw_payload_qos,
    output wire [31:0] M_AXI_GP0_w_payload_data,
    output wire [3:0] M_AXI_GP0_w_payload_strb,
    output wire M_AXI_GP0_w_payload_last,
    input wire [11:0] M_AXI_GP0_r_payload_id,
    input wire M_AXI_GP0_r_payload_last,
    input wire [1:0] M_AXI_GP0_r_payload_resp,
    input wire [31:0] M_AXI_GP0_r_payload_data,
    input wire [11:0] M_AXI_GP0_b_payload_id,
    input wire [1:0] M_AXI_GP0_b_payload_resp,
  `endif
  `ifdef PS_MASTER_AXI_GP1
    //M_AXI_GP1
    output wire M_AXI_GP1_ARESET,
    output wire M_AXI_GP1_ARVALID,
    output wire M_AXI_GP1_AWVALID,
    output wire M_AXI_GP1_BREADY,
    output wire M_AXI_GP1_RREADY,
    output wire M_AXI_GP1_WLAST,
    output wire M_AXI_GP1_WVALID,
    output wire [11:0] M_AXI_GP1_ARID,
    output wire [11:0] M_AXI_GP1_AWID,
    output wire [11:0] M_AXI_GP1_WID,
    output wire [1:0] M_AXI_GP1_ARBURST,
    output wire [1:0] M_AXI_GP1_ARLOCK,
    output wire [1:0] M_AXI_GP1_ARSIZE,
    output wire [1:0] M_AXI_GP1_AWBURST,
    output wire [1:0] M_AXI_GP1_AWLOCK,
    output wire [1:0] M_AXI_GP1_AWSIZE,
    output wire [2:0] M_AXI_GP1_ARPROT,
    output wire [2:0] M_AXI_GP1_AWPROT,
    output wire [31:0] M_AXI_GP1_ARADDR,
    output wire [31:0] M_AXI_GP1_AWADDR,
    output wire [31:0] M_AXI_GP1_WDATA,
    output wire [3:0] M_AXI_GP1_ARCACHE,
    output wire [3:0] M_AXI_GP1_ARLEN,
    output wire [3:0] M_AXI_GP1_ARQOS,
    output wire [3:0] M_AXI_GP1_AWCACHE,
    output wire [3:0] M_AXI_GP1_AWLEN,
    output wire [3:0] M_AXI_GP1_AWQOS,
    output wire [3:0] M_AXI_GP1_WSTRB,
    input wire M_AXI_GP1_ACLK,
    input wire M_AXI_GP1_ARREADY,
    input wire M_AXI_GP1_AWREADY,
    input wire M_AXI_GP1_BVALID,
    input wire M_AXI_GP1_RLAST,
    input wire M_AXI_GP1_RVALID,
    input wire M_AXI_GP1_WREADY,  
    input wire [11:0] M_AXI_GP1_BID,
    input wire [11:0] M_AXI_GP1_RID,
    input wire [1:0] M_AXI_GP1_BRESP,
    input wire [1:0] M_AXI_GP1_RRESP,
    input wire [31:0] M_AXI_GP1_RDATA,
  `endif
  `ifdef PS_SLAVE_AXI_GP0
    // S_AXI_GP0
    output wire S_AXI_GP0_ARESET,
    output wire S_AXI_GP0_ARREADY,
    output wire S_AXI_GP0_AWREADY,
    output wire S_AXI_GP0_BVALID,
    output wire S_AXI_GP0_RLAST,
    output wire S_AXI_GP0_RVALID,
    output wire S_AXI_GP0_WREADY,  
    output wire [1:0] S_AXI_GP0_BRESP,
    output wire [1:0] S_AXI_GP0_RRESP,
    output wire [31:0] S_AXI_GP0_RDATA,
    output wire [5:0] S_AXI_GP0_BID,
    output wire [5:0] S_AXI_GP0_RID,
    input wire S_AXI_GP0_ACLK,
    input wire S_AXI_GP0_ARVALID,
    input wire S_AXI_GP0_AWVALID,
    input wire S_AXI_GP0_BREADY,
    input wire S_AXI_GP0_RREADY,
    input wire S_AXI_GP0_WLAST,
    input wire S_AXI_GP0_WVALID,
    input wire [1:0] S_AXI_GP0_ARBURST,
    input wire [1:0] S_AXI_GP0_ARLOCK,
    input wire [1:0] S_AXI_GP0_ARSIZE,
    input wire [1:0] S_AXI_GP0_AWBURST,
    input wire [1:0] S_AXI_GP0_AWLOCK,
    input wire [1:0] S_AXI_GP0_AWSIZE,
    input wire [2:0] S_AXI_GP0_ARPROT,
    input wire [2:0] S_AXI_GP0_AWPROT,
    input wire [31:0] S_AXI_GP0_ARADDR,
    input wire [31:0] S_AXI_GP0_AWADDR,
    input wire [31:0] S_AXI_GP0_WDATA,
    input wire [3:0] S_AXI_GP0_ARCACHE,
    input wire [3:0] S_AXI_GP0_ARLEN,
    input wire [3:0] S_AXI_GP0_ARQOS,
    input wire [3:0] S_AXI_GP0_AWCACHE,
    input wire [3:0] S_AXI_GP0_AWLEN,
    input wire [3:0] S_AXI_GP0_AWQOS,
    input wire [3:0] S_AXI_GP0_WSTRB,
    input wire [5:0] S_AXI_GP0_ARID,
    input wire [5:0] S_AXI_GP0_AWID,
    input wire [5:0] S_AXI_GP0_WID,  
  `endif
  `ifdef PS_SLAVE_AXI_GP1
    // S_AXI_GP1
    output wire S_AXI_GP1_ARESET,
    output wire S_AXI_GP1_ARREADY,
    output wire S_AXI_GP1_AWREADY,
    output wire S_AXI_GP1_BVALID,
    output wire S_AXI_GP1_RLAST,
    output wire S_AXI_GP1_RVALID,
    output wire S_AXI_GP1_WREADY,  
    output wire [1:0] S_AXI_GP1_BRESP,
    output wire [1:0] S_AXI_GP1_RRESP,
    output wire [31:0] S_AXI_GP1_RDATA,
    output wire [5:0] S_AXI_GP1_BID,
    output wire [5:0] S_AXI_GP1_RID,
    input wire S_AXI_GP1_ACLK,
    input wire S_AXI_GP1_ARVALID,
    input wire S_AXI_GP1_AWVALID,
    input wire S_AXI_GP1_BREADY,
    input wire S_AXI_GP1_RREADY,
    input wire S_AXI_GP1_WLAST,
    input wire S_AXI_GP1_WVALID,
    input wire [1:0] S_AXI_GP1_ARBURST,
    input wire [1:0] S_AXI_GP1_ARLOCK,
    input wire [1:0] S_AXI_GP1_ARSIZE,
    input wire [1:0] S_AXI_GP1_AWBURST,
    input wire [1:0] S_AXI_GP1_AWLOCK,
    input wire [1:0] S_AXI_GP1_AWSIZE,
    input wire [2:0] S_AXI_GP1_ARPROT,
    input wire [2:0] S_AXI_GP1_AWPROT,
    input wire [31:0] S_AXI_GP1_ARADDR,
    input wire [31:0] S_AXI_GP1_AWADDR,
    input wire [31:0] S_AXI_GP1_WDATA,
    input wire [3:0] S_AXI_GP1_ARCACHE,
    input wire [3:0] S_AXI_GP1_ARLEN,
    input wire [3:0] S_AXI_GP1_ARQOS,
    input wire [3:0] S_AXI_GP1_AWCACHE,
    input wire [3:0] S_AXI_GP1_AWLEN,
    input wire [3:0] S_AXI_GP1_AWQOS,
    input wire [3:0] S_AXI_GP1_WSTRB,
    input wire [5:0] S_AXI_GP1_ARID,
    input wire [5:0] S_AXI_GP1_AWID,
    input wire [5:0] S_AXI_GP1_WID, 
  `endif
  `ifdef PS_SLAVE_AXI_ACP
    //S_AXI_ACP
    output wire S_AXI_ACP_ARESET,
    output wire S_AXI_ACP_ARREADY,
    output wire S_AXI_ACP_AWREADY,
    output wire S_AXI_ACP_BVALID,
    output wire S_AXI_ACP_RLAST,
    output wire S_AXI_ACP_RVALID,
    output wire S_AXI_ACP_WREADY,  
    output wire [1:0] S_AXI_ACP_BRESP,
    output wire [1:0] S_AXI_ACP_RRESP,
    output wire [2 : 0] S_AXI_ACP_BID,
    output wire [2 : 0] S_AXI_ACP_RID,
    output wire [63:0] S_AXI_ACP_RDATA,
    input wire S_AXI_ACP_ACLK,
    input wire S_AXI_ACP_ARVALID,
    input wire S_AXI_ACP_AWVALID,
    input wire S_AXI_ACP_BREADY,
    input wire S_AXI_ACP_RREADY,
    input wire S_AXI_ACP_WLAST,
    input wire S_AXI_ACP_WVALID,
    input wire [2:0] S_AXI_ACP_ARID,
    input wire [2:0] S_AXI_ACP_ARPROT,
    input wire [2:0] S_AXI_ACP_AWID,
    input wire [2:0] S_AXI_ACP_AWPROT,
    input wire [2:0] S_AXI_ACP_WID,
    input wire [31:0] S_AXI_ACP_ARADDR,
    input wire [31:0] S_AXI_ACP_AWADDR,
    input wire [3:0] S_AXI_ACP_ARCACHE,
    input wire [3:0] S_AXI_ACP_ARLEN,
    input wire [3:0] S_AXI_ACP_ARQOS,
    input wire [3:0] S_AXI_ACP_AWCACHE,
    input wire [3:0] S_AXI_ACP_AWLEN,
    input wire [3:0] S_AXI_ACP_AWQOS,
    input wire [1:0] S_AXI_ACP_ARBURST,
    input wire [1:0] S_AXI_ACP_ARLOCK,
    input wire [1:0] S_AXI_ACP_ARSIZE,
    input wire [1:0] S_AXI_ACP_AWBURST,
    input wire [1:0] S_AXI_ACP_AWLOCK,
    input wire [1:0] S_AXI_ACP_AWSIZE,
    input wire [4:0] S_AXI_ACP_ARUSER,
    input wire [4:0] S_AXI_ACP_AWUSER,
    input wire [63:0] S_AXI_ACP_WDATA,
    input wire [7:0] S_AXI_ACP_WSTRB, 
  `endif
  `ifdef PS_SLAVE_AXI_HP0
    // AXI HP0
    output wire S_AXI_HP0_ARESET,
    output wire S_AXI_HP0_ARREADY,
    output wire S_AXI_HP0_AWREADY,
    output wire S_AXI_HP0_BVALID,
    output wire S_AXI_HP0_RLAST,
    output wire S_AXI_HP0_RVALID,
    output wire S_AXI_HP0_WREADY,  
    output wire [1:0] S_AXI_HP0_BRESP,
    output wire [1:0] S_AXI_HP0_RRESP,
    output wire [5:0] S_AXI_HP0_BID,
    output wire [5:0] S_AXI_HP0_RID,
    output wire [63:0] S_AXI_HP0_RDATA,
    output wire [7:0] S_AXI_HP0_RCOUNT,
    output wire [7:0] S_AXI_HP0_WCOUNT,
    output wire [2:0] S_AXI_HP0_RACOUNT,
    output wire [5:0] S_AXI_HP0_WACOUNT,
    input wire S_AXI_HP0_ACLK,
    input wire S_AXI_HP0_ARVALID,
    input wire S_AXI_HP0_AWVALID,
    input wire S_AXI_HP0_BREADY,
    input wire S_AXI_HP0_RDISSUECAP1_EN,
    input wire S_AXI_HP0_RREADY,
    input wire S_AXI_HP0_WLAST,
    input wire S_AXI_HP0_WRISSUECAP1_EN,
    input wire S_AXI_HP0_WVALID,
    input wire [1:0] S_AXI_HP0_ARBURST,
    input wire [1:0] S_AXI_HP0_ARLOCK,
    input wire [1:0] S_AXI_HP0_ARSIZE,
    input wire [1:0] S_AXI_HP0_AWBURST,
    input wire [1:0] S_AXI_HP0_AWLOCK,
    input wire [1:0] S_AXI_HP0_AWSIZE,
    input wire [2:0] S_AXI_HP0_ARPROT,
    input wire [2:0] S_AXI_HP0_AWPROT,
    input wire [31:0] S_AXI_HP0_ARADDR,
    input wire [31:0] S_AXI_HP0_AWADDR,
    input wire [3:0] S_AXI_HP0_ARCACHE,
    input wire [3:0] S_AXI_HP0_ARLEN,
    input wire [3:0] S_AXI_HP0_ARQOS,
    input wire [3:0] S_AXI_HP0_AWCACHE,
    input wire [3:0] S_AXI_HP0_AWLEN,
    input wire [3:0] S_AXI_HP0_AWQOS,
    input wire [5:0] S_AXI_HP0_ARID,
    input wire [5:0] S_AXI_HP0_AWID,
    input wire [5:0] S_AXI_HP0_WID,
    input wire [63:0] S_AXI_HP0_WDATA,
    input wire [7:0] S_AXI_HP0_WSTRB,
  `endif
  `ifdef PS_SLAVE_AXI_HP1
    // AXI HP1
    output wire S_AXI_HP1_ARESET,
    output wire S_AXI_HP1_ARREADY,
    output wire S_AXI_HP1_AWREADY,
    output wire S_AXI_HP1_BVALID,
    output wire S_AXI_HP1_RLAST,
    output wire S_AXI_HP1_RVALID,
    output wire S_AXI_HP1_WREADY,  
    output wire [1:0] S_AXI_HP1_BRESP,
    output wire [1:0] S_AXI_HP1_RRESP,
    output wire [5:0] S_AXI_HP1_BID,
    output wire [5:0] S_AXI_HP1_RID,
    output wire [63:0] S_AXI_HP1_RDATA,
    output wire [7:0] S_AXI_HP1_RCOUNT,
    output wire [7:0] S_AXI_HP1_WCOUNT,
    output wire [2:0] S_AXI_HP1_RACOUNT,
    output wire [5:0] S_AXI_HP1_WACOUNT,
    input wire S_AXI_HP1_ACLK,
    input wire S_AXI_HP1_ARVALID,
    input wire S_AXI_HP1_AWVALID,
    input wire S_AXI_HP1_BREADY,
    input wire S_AXI_HP1_RDISSUECAP1_EN,
    input wire S_AXI_HP1_RREADY,
    input wire S_AXI_HP1_WLAST,
    input wire S_AXI_HP1_WRISSUECAP1_EN,
    input wire S_AXI_HP1_WVALID,
    input wire [1:0] S_AXI_HP1_ARBURST,
    input wire [1:0] S_AXI_HP1_ARLOCK,
    input wire [1:0] S_AXI_HP1_ARSIZE,
    input wire [1:0] S_AXI_HP1_AWBURST,
    input wire [1:0] S_AXI_HP1_AWLOCK,
    input wire [1:0] S_AXI_HP1_AWSIZE,
    input wire [2:0] S_AXI_HP1_ARPROT,
    input wire [2:0] S_AXI_HP1_AWPROT,
    input wire [31:0] S_AXI_HP1_ARADDR,
    input wire [31:0] S_AXI_HP1_AWADDR,
    input wire [3:0] S_AXI_HP1_ARCACHE,
    input wire [3:0] S_AXI_HP1_ARLEN,
    input wire [3:0] S_AXI_HP1_ARQOS,
    input wire [3:0] S_AXI_HP1_AWCACHE,
    input wire [3:0] S_AXI_HP1_AWLEN,
    input wire [3:0] S_AXI_HP1_AWQOS,
    input wire [5:0] S_AXI_HP1_ARID,
    input wire [5:0] S_AXI_HP1_AWID,
    input wire [5:0] S_AXI_HP1_WID,
    input wire [63:0] S_AXI_HP1_WDATA,
    input wire [7:0] S_AXI_HP1_WSTRB,
  `endif
  `ifdef PS_SLAVE_AXI_HP2
    // S_AXI_HP2
    output wire S_AXI_HP2_ARESET,
    output wire S_AXI_HP2_ARREADY,
    output wire S_AXI_HP2_AWREADY,
    output wire S_AXI_HP2_BVALID,
    output wire S_AXI_HP2_RLAST,
    output wire S_AXI_HP2_RVALID,
    output wire S_AXI_HP2_WREADY,  
    output wire [1:0] S_AXI_HP2_BRESP,
    output wire [1:0] S_AXI_HP2_RRESP,
    output wire [5:0] S_AXI_HP2_BID,
    output wire [5:0] S_AXI_HP2_RID,
    output wire [63:0] S_AXI_HP2_RDATA,
    output wire [7:0] S_AXI_HP2_RCOUNT,
    output wire [7:0] S_AXI_HP2_WCOUNT,
    output wire [2:0] S_AXI_HP2_RACOUNT,
    output wire [5:0] S_AXI_HP2_WACOUNT,
    input wire S_AXI_HP2_ACLK,
    input wire S_AXI_HP2_ARVALID,
    input wire S_AXI_HP2_AWVALID,
    input wire S_AXI_HP2_BREADY,
    input wire S_AXI_HP2_RDISSUECAP1_EN,
    input wire S_AXI_HP2_RREADY,
    input wire S_AXI_HP2_WLAST,
    input wire S_AXI_HP2_WRISSUECAP1_EN,
    input wire S_AXI_HP2_WVALID,
    input wire [1:0] S_AXI_HP2_ARBURST,
    input wire [1:0] S_AXI_HP2_ARLOCK,
    input wire [1:0] S_AXI_HP2_ARSIZE,
    input wire [1:0] S_AXI_HP2_AWBURST,
    input wire [1:0] S_AXI_HP2_AWLOCK,
    input wire [1:0] S_AXI_HP2_AWSIZE,
    input wire [2:0] S_AXI_HP2_ARPROT,
    input wire [2:0] S_AXI_HP2_AWPROT,
    input wire [31:0] S_AXI_HP2_ARADDR,
    input wire [31:0] S_AXI_HP2_AWADDR,
    input wire [3:0] S_AXI_HP2_ARCACHE,
    input wire [3:0] S_AXI_HP2_ARLEN,
    input wire [3:0] S_AXI_HP2_ARQOS,
    input wire [3:0] S_AXI_HP2_AWCACHE,
    input wire [3:0] S_AXI_HP2_AWLEN,
    input wire [3:0] S_AXI_HP2_AWQOS,
    input wire [5:0] S_AXI_HP2_ARID,
    input wire [5:0] S_AXI_HP2_AWID,
    input wire [5:0] S_AXI_HP2_WID,
    input wire [63:0] S_AXI_HP2_WDATA,
    input wire [7:0] S_AXI_HP2_WSTRB,
  `endif
  `ifdef PS_SLAVE_AXI_HP3
    // S_AXI_HP_3
    output wire S_AXI_HP3_ARESET,
    output wire S_AXI_HP3_ARREADY,
    output wire S_AXI_HP3_AWREADY,
    output wire S_AXI_HP3_BVALID,
    output wire S_AXI_HP3_RLAST,
    output wire S_AXI_HP3_RVALID,
    output wire S_AXI_HP3_WREADY,  
    output wire [1:0] S_AXI_HP3_BRESP,
    output wire [1:0] S_AXI_HP3_RRESP,
    output wire [5:0] S_AXI_HP3_BID,
    output wire [5:0] S_AXI_HP3_RID,
    output wire [63:0] S_AXI_HP3_RDATA,
    output wire [7:0] S_AXI_HP3_RCOUNT,
    output wire [7:0] S_AXI_HP3_WCOUNT,
    output wire [2:0] S_AXI_HP3_RACOUNT,
    output wire [5:0] S_AXI_HP3_WACOUNT,
    input wire S_AXI_HP3_ACLK,
    input wire S_AXI_HP3_ARVALID,
    input wire S_AXI_HP3_AWVALID,
    input wire S_AXI_HP3_BREADY,
    input wire S_AXI_HP3_RDISSUECAP1_EN,
    input wire S_AXI_HP3_RREADY,
    input wire S_AXI_HP3_WLAST,
    input wire S_AXI_HP3_WRISSUECAP1_EN,
    input wire S_AXI_HP3_WVALID,
    input wire [1:0] S_AXI_HP3_ARBURST,
    input wire [1:0] S_AXI_HP3_ARLOCK,
    input wire [1:0] S_AXI_HP3_ARSIZE,
    input wire [1:0] S_AXI_HP3_AWBURST,
    input wire [1:0] S_AXI_HP3_AWLOCK,
    input wire [1:0] S_AXI_HP3_AWSIZE,
    input wire [2:0] S_AXI_HP3_ARPROT,
    input wire [2:0] S_AXI_HP3_AWPROT,
    input wire [31:0] S_AXI_HP3_ARADDR,
    input wire [31:0] S_AXI_HP3_AWADDR,
    input wire [3:0] S_AXI_HP3_ARCACHE,
    input wire [3:0] S_AXI_HP3_ARLEN,
    input wire [3:0] S_AXI_HP3_ARQOS,
    input wire [3:0] S_AXI_HP3_AWCACHE,
    input wire [3:0] S_AXI_HP3_AWLEN,
    input wire [3:0] S_AXI_HP3_AWQOS,
    input wire [5:0] S_AXI_HP3_ARID,
    input wire [5:0] S_AXI_HP3_AWID,
    input wire [5:0] S_AXI_HP3_WID,
    input wire [63:0] S_AXI_HP3_WDATA,
    input wire [7:0] S_AXI_HP3_WSTRB,
  `endif
  // DDR
  input [3:0] DDR_ARB,
  inout wire DDR_CAS_n,
  inout wire DDR_CKE,
  inout wire DDR_Clk_n,
  inout wire DDR_Clk,
  inout wire DDR_CS_n,
  inout wire DDR_DRSTB,
  inout wire DDR_ODT,
  inout wire DDR_RAS_n,
  inout wire DDR_WEB,
  inout wire [2:0]  DDR_BankAddr,
  inout wire [14:0] DDR_Addr,
  inout wire DDR_VRN,
  inout wire DDR_VRP,
  inout wire [3:0]  DDR_DM,
  inout wire [31:0] DDR_DQ,
  inout wire [3:0]  DDR_DQS_n,
  inout wire [3:0]  DDR_DQS,

  // PS Clock and Reset wires
  output wire PS_SYSTEM_RESET,
  output wire PS_CLK,         
  output wire PS_POWER_ON_RESET
  
);
  `ifdef PS_MASTER_AXI_GP0
    wire [1:0] M_AXI_GP0_ar_payload_lock_adaptor; // Axi4 lock simplified
    wire [1:0] M_AXI_GP0_aw_payload_lock_adaptor;
    wire [1:0] M_AXI_GP0_ar_payload_size_adaptor; // size can't be larger than bus so pad with 0
    wire [1:0] M_AXI_GP0_aw_payload_size_adaptor;
    wire [3:0] M_AXI_GP0_ar_payload_len_adaptor; // axi4 can issue longer burst we don't so pad with 0
    wire [3:0] M_AXI_GP0_aw_payload_len_adaptor;

    wire [11:0] M_AXI_GP0_w_payload_id; // not used for Axi4
    assign M_AXI_GP0_ar_payload_lock = M_AXI_GP0_ar_payload_lock_adaptor[0];
    assign M_AXI_GP0_aw_payload_lock = M_AXI_GP0_aw_payload_lock_adaptor[0];
    assign M_AXI_GP0_ar_payload_size = { 1'b0, M_AXI_GP0_ar_payload_size_adaptor };
    assign M_AXI_GP0_aw_payload_size = { 1'b0, M_AXI_GP0_aw_payload_size_adaptor };
    assign M_AXI_GP0_ar_payload_len = { 4'h0, M_AXI_GP0_ar_payload_len_adaptor };
    assign M_AXI_GP0_aw_payload_len = { 4'h0, M_AXI_GP0_aw_payload_len_adaptor };      
  `endif

  // ----- Instaniate the PS7 wrapper
  ps7_wrapper ps7_wrapper_i (
  `ifdef USE_CAN0
    .CAN0_PHY_TX(CAN0_PHY_TX),
    .CAN0_PHY_RX(CAN0_PHY_RX),
  `endif

  `ifdef USE_CAN1
    .CAN1_PHY_TX(CAN1_PHY_TX),
    .CAN1_PHY_RX(CAN1_PHY_RX),
  `endif

  `ifdef USE_ENET0
    .ENET0_GMII_TX_EN(ENET0_GMII_TX_EN_i),
    .ENET0_GMII_TX_ER(ENET0_GMII_TX_ER_i),
    .ENET0_GMII_RX_CLK(ENET0_GMII_RX_CLK),
    .ENET0_GMII_TX_CLK(ENET0_GMII_TX_CLK),
    .ENET0_GMII_TXD(ENET0_GMII_TXD_i),
    .ENET0_GMII_COL(ENET0_GMII_COL_o),
    .ENET0_GMII_CRS(ENET0_GMII_CRS_o),
    .ENET0_GMII_RX_DV(ENET0_GMII_RX_DV_o),
    .ENET0_GMII_RX_ER(ENET0_GMII_RX_ER_o),
    .ENET0_GMII_RXD(ENET0_GMII_RXD_o),
    .ENET0_MDIO_MDC(ENET0_MDIO_MDC),
    .ENET0_MDIO_O(ENET0_MDIO_O),
    .ENET0_MDIO_T_n(ENET0_MDIO_T_n),
    .ENET0_PTP_DELAY_REQ_RX(ENET0_PTP_DELAY_REQ_RX),
    .ENET0_PTP_DELAY_REQ_TX(ENET0_PTP_DELAY_REQ_TX),
    .ENET0_PTP_PDELAY_REQ_RX(ENET0_PTP_PDELAY_REQ_RX),
    .ENET0_PTP_PDELAY_REQ_TX(ENET0_PTP_PDELAY_REQ_TX),
    .ENET0_PTP_PDELAY_RESP_RX(ENET0_PTP_PDELAY_RESP_RX),
    .ENET0_PTP_PDELAY_RESP_TX(ENET0_PTP_PDELAY_RESP_TX),
    .ENET0_PTP_SYNC_FRAME_RX(ENET0_PTP_SYNC_FRAME_RX),
    .ENET0_PTP_SYNC_FRAME_TX(ENET0_PTP_SYNC_FRAME_TX),
    .ENET0_SOF_RX(ENET0_SOF_RX),
    .ENET0_SOF_TX(ENET0_SOF_TX),
    .ENET0_MDIO_I(ENET0_MDIO_I),
    .ENET0_EXT_INTIN(ENET0_EXT_INTIN),
  `endif
  `ifdef USE_ENET1
    .ENET1_GMII_TX_EN(ENET1_GMII_TX_EN_i),
    .ENET1_GMII_TX_ER(ENET1_GMII_TX_ER_i),
    .ENET1_GMII_RX_CLK(ENET1_GMII_RX_CLK),
    .ENET1_GMII_TX_CLK(ENET1_GMII_TX_CLK),
    .ENET1_GMII_TXD(ENET1_GMII_TXD_i),
    .ENET1_GMII_COL(ENET1_GMII_COL_o),
    .ENET1_GMII_CRS(ENET1_GMII_CRS_o),
    .ENET1_GMII_RX_DV(ENET1_GMII_RX_DV_o),
    .ENET1_GMII_RX_ER(ENET1_GMII_RX_ER_o),
    .ENET1_GMII_RXD(ENET1_GMII_RXD_o),
    .ENET1_MDIO_MDC(ENET1_MDIO_MDC),
    .ENET1_MDIO_O(ENET1_MDIO_O),
    .ENET1_MDIO_T_n(ENET1_MDIO_T_n),
    .ENET1_PTP_DELAY_REQ_RX(ENET1_PTP_DELAY_REQ_RX),
    .ENET1_PTP_DELAY_REQ_TX(ENET1_PTP_DELAY_REQ_TX),
    .ENET1_PTP_PDELAY_REQ_RX(ENET1_PTP_PDELAY_REQ_RX),
    .ENET1_PTP_PDELAY_REQ_TX(ENET1_PTP_PDELAY_REQ_TX),
    .ENET1_PTP_PDELAY_RESP_RX(ENET1_PTP_PDELAY_RESP_RX),
    .ENET1_PTP_PDELAY_RESP_TX(ENET1_PTP_PDELAY_RESP_TX),
    .ENET1_PTP_SYNC_FRAME_RX(ENET1_PTP_SYNC_FRAME_RX),
    .ENET1_PTP_SYNC_FRAME_TX(ENET1_PTP_SYNC_FRAME_TX),
    .ENET1_SOF_RX(ENET1_SOF_RX),
    .ENET1_SOF_TX(ENET1_SOF_TX),
    .ENET1_MDIO_I(ENET1_MDIO_I),
    .ENET1_EXT_INTIN(ENET1_EXT_INTIN),
  `endif
  `ifdef USE_DMA0
	  .DMA0_ACLK		            (DMA0_ACLK),
	  .DMA0_RESET_n		          (DMA0_RESET_n),  
	  .DMA0_DATYPE		          (DMA0_DATYPE),
	  .DMA0_DAVALID		          (DMA0_DAVALID),
	  .DMA0_DRREADY		          (DMA0_DRREADY),  
	  .DMA0_DAREADY		          (DMA0_DAREADY),
	  .DMA0_DRLAST		          (DMA0_DRLAST),
	  .DMA0_DRTYPE              (DMA0_DRTYPE),
	  .DMA0_DRVALID		          (DMA0_DRVALID),
  `endif
  `ifdef USE_DMA1
	  .DMA1_ACLK		            (DMA1_ACLK),
	  .DMA1_RESET_n		          (DMA1_RESET_n),
	  .DMA1_DATYPE		          (DMA1_DATYPE),
	  .DMA1_DAVALID		          (DMA1_DAVALID),
	  .DMA1_DRREADY		          (DMA1_DRREADY),
	  .DMA1_DAREADY		          (DMA1_DAREADY),
	  .DMA1_DRLAST		          (DMA1_DRLAST),
	  .DMA1_DRTYPE              (DMA1_DRTYPE),  
	  .DMA1_DRVALID		          (DMA1_DRVALID),
  `endif
  `ifdef USE_DMA2
	  .DMA2_ACLK		            (DMA2_ACLK),
	  .DMA2_RESET_n		          (DMA2_RESET_n),
	  .DMA2_DATYPE		          (DMA2_DATYPE),
	  .DMA2_DAVALID		          (DMA2_DAVALID),
	  .DMA2_DRREADY		          (DMA2_DRREADY),
	  .DMA2_DAREADY		          (DMA2_DAREADY),
	  .DMA2_DRLAST		          (DMA2_DRLAST),
	  .DMA2_DRTYPE              (DMA2_DRTYPE),    
	  .DMA2_DRVALID		          (DMA2_DRVALID),
  `endif
  `ifdef USE_DMA3
	  .DMA3_ACLK		            (DMA3_ACLK),
	  .DMA3_RESET_n		          (DMA3_RESET_n),
	  .DMA3_DAREADY		          (DMA3_DAREADY),
	  .DMA3_DRLAST		          (DMA3_DRLAST),
	  .DMA3_DRTYPE              (DMA3_DRTYPE),
	  .DMA3_DRVALID		          (DMA3_DRVALID),
	  .DMA3_DATYPE		          (DMA3_DATYPE),
	  .DMA3_DAVALID		          (DMA3_DAVALID),
	  .DMA3_DRREADY		          (DMA3_DRREADY),
  `endif
  `ifdef USE_GPIO
    .GPIO_I                   (GPIO_I),
    .GPIO_O                   (GPIO_O),
    .GPIO_T_n                 (GPIO_T_n),
  `endif
  `ifdef USE_MIO
    .MIO                      (MIO),
  `endif

  `ifdef USE_I2C0
    .I2C0_SDA_I               (I2C0_SDA_I),
    .I2C0_SDA_O               (I2C0_SDA_O),
    .I2C0_SDA_T               (I2C0_SDA_T),
    .I2C0_SCL_I               (I2C0_SCL_I),
    .I2C0_SCL_O               (I2C0_SCL_O),
    .I2C0_SCL_T               (I2C0_SCL_T),
  `endif    
  `ifdef USE_I2C1
    .I2C1_SDA_I               (I2C1_SDA_I),
    .I2C1_SDA_O               (I2C1_SDA_O),
    .I2C1_SDA_T               (I2C1_SDA_T),
    .I2C1_SCL_I               (I2C1_SCL_I),
    .I2C1_SCL_O               (I2C1_SCL_O),
    .I2C1_SCL_T               (I2C1_SCL_T),
  `endif
  `ifdef USE_SDIO0
    .SDIO0_CLK                (SDIO0_CLK),
    .SDIO0_CLK_FB             (SDIO0_CLK_FB),
    .SDIO0_CMD_O              (SDIO0_CMD_O),
    .SDIO0_CMD_I              (SDIO0_CMD_I),
    .SDIO0_CMD_T              (SDIO0_CMD_T),
    .SDIO0_DATA_I             (SDIO0_DATA_I),
    .SDIO0_DATA_O             (SDIO0_DATA_O),
    .SDIO0_DATA_T             (SDIO0_DATA_T),
    .SDIO0_LED                (SDIO0_LED),
    .SDIO0_CDN                (SDIO0_CDN),
    .SDIO0_WP                 (SDIO0_WP),  
    .SDIO0_BUSPOW             (SDIO0_BUSPOW),
    .SDIO0_BUSVOLT            (SDIO0_BUSVOLT),
  `endif
  `ifdef USE_SDIO1
    .SDIO1_CLK                (SDIO1_CLK),
    .SDIO1_CLK_FB             (SDIO1_CLK_FB),
    .SDIO1_CMD_O              (SDIO1_CMD_O),
    .SDIO1_CMD_I              (SDIO1_CMD_I),
    .SDIO1_CMD_T              (SDIO1_CMD_T),
    .SDIO1_DATA_I             (SDIO1_DATA_I),
    .SDIO1_DATA_O             (SDIO1_DATA_O),
    .SDIO1_DATA_T             (SDIO1_DATA_T),
    .SDIO1_LED                (SDIO1_LED),
    .SDIO1_CDN                (SDIO1_CDN),
    .SDIO1_WP                 (SDIO1_WP),
    .SDIO1_BUSPOW             (SDIO1_BUSPOW),
    .SDIO1_BUSVOLT            (SDIO1_BUSVOLT),
  `endif
  `ifdef USE_SPI0
      // SPI wires
    .SPI0_SCLK_I              (SPI0_SCLK_I),
    .SPI0_SCLK_O              (SPI0_SCLK_O),
    .SPI0_SCLK_T              (SPI0_SCLK_T_n),
    .SPI0_MOSI_I              (SPI0_MOSI_I),
    .SPI0_MOSI_O              (SPI0_MOSI_O),
    .SPI0_MOSI_T              (SPI0_MOSI_T),
    .SPI0_MISO_I              (SPI0_MISO_I),
    .SPI0_MISO_O              (SPI0_MISO_O),
    .SPI0_MISO_T              (SPI0_MISO_T),
    .SPI0_SS_I                (SPI0_SS_I),
    .SPI0_SS_O                (SPI0_SS_O),
    .SPI0_SS1_O               (SPI0_SS1_O),
    .SPI0_SS2_O               (SPI0_SS2_O),
    .SPI0_SS_T                (SPI0_SS_T),
  `endif
  `ifdef USE_SPI1
    .SPI1_SCLK_I              (SPI1_SCLK_I),
    .SPI1_SCLK_O              (SPI1_SCLK_O),
    .SPI1_SCLK_T              (SPI1_SCLK_T),
    .SPI1_MOSI_I              (SPI1_MOSI_I),
    .SPI1_MOSI_O              (SPI1_MOSI_O),
    .SPI1_MOSI_T              (SPI1_MOSI_T),
    .SPI1_MISO_I              (SPI1_MISO_I),
    .SPI1_MISO_O              (SPI1_MISO_O),
    .SPI1_MISO_T              (SPI1_MISO_T),
    .SPI1_SS_I                (SPI1_SS_I),
    .SPI1_SS_O                (SPI1_SS_O),
    .SPI1_SS1_O               (SPI1_SS1_O),
    .SPI1_SS2_O               (SPI1_SS2_O),
    .SPI1_SS_T                (SPI1_SS_T),
  `endif
  `ifdef USE_UART0
    .UART0_DTRN               (UART0_DTRN),
    .UART0_RTSN               (UART0_RTSN), 
    .UART0_TX                 (UART0_TX),
    .UART0_CTSN               (UART0_CTSN),
    .UART0_DCDN               (UART0_DCDN),
    .UART0_DSRN               (UART0_DSRN),
    .UART0_RIN                (UART0_RIN),
    .UART0_RX                 (UART0_RX),
  `endif
  `ifdef USE_UART1
    .UART1_DTRN               (UART1_DTRN),
    .UART1_RX                 (UART1_RX),
    .UART1_RTSN               (UART1_RTSN),  
    .UART1_TX                 (UART1_TX),
    .UART1_CTSN               (UART1_CTSN),
    .UART1_DCDN               (UART1_DCDN),
    .UART1_DSRN               (UART1_DSRN),
    .UART1_RIN                (UART1_RIN),
  `endif
  `ifdef USE_JTAG
    .PJTAG_TCK                (PJTAG_TCK),
    .PJTAG_TMS                (PJTAG_TMS),
    .PJTAG_TDI                (PJTAG_TDI),
    .PJTAG_TDO_O              (PJTAG_TDO_O),
    .PJTAG_TDO_T              (PJTAG_TDO_T),
  `endif
  `ifdef USE_TTC0
    .TTC0_WAVE0_OUT           (TTC0_WAVE0_OUT),
    .TTC0_WAVE1_OUT           (TTC0_WAVE1_OUT),
    .TTC0_WAVE2_OUT           (TTC0_WAVE2_OUT),
    .TTC0_CLK0_IN             (TTC0_CLK0_IN),
    .TTC0_CLK1_IN             (TTC0_CLK1_IN),
    .TTC0_CLK2_IN             (TTC0_CLK2_IN),
  `endif
  `ifdef USE_TTC1
    .TTC1_WAVE0_OUT           (TTC1_WAVE0_OUT),
    .TTC1_WAVE1_OUT           (TTC1_WAVE1_OUT),
    .TTC1_WAVE2_OUT           (TTC1_WAVE2_OUT),
    .TTC1_CLK0_IN             (TTC1_CLK0_IN),
    .TTC1_CLK1_IN             (TTC1_CLK1_IN),
    .TTC1_CLK2_IN             (TTC1_CLK2_IN),
  `endif
  `ifdef USE_TRACE
    .TRACE_CLK                (TRACE_CLK),
    .TRACE_CTL                (TRACE_CTL),
    .TRACE_DATA               (TRACE_DATA),
    .TRACE_CLK_OUT            (TRACE_CLK_OUT),
    .FTMD_TRACEIN_DATA        (FTMD_TRACEIN_DATA),
    .FTMD_TRACEIN_VALID       (FTMD_TRACEIN_VALID),
    .FTMD_TRACEIN_CLK         (FTMD_TRACEIN_CLK),
    .FTMD_TRACEIN_ATID        (FTMD_TRACEIN_ATID),
    .FTMT_F2P_TRIG_0          (FTMT_F2P_TRIG_0),
    .FTMT_F2P_TRIGACK_0       (FTMT_F2P_TRIGACK_0),
    .FTMT_F2P_TRIG_1          (FTMT_F2P_TRIG_1),
    .FTMT_F2P_TRIGACK_1       (FTMT_F2P_TRIGACK_1),
    .FTMT_F2P_TRIG_2          (FTMT_F2P_TRIG_2),
    .FTMT_F2P_TRIGACK_2       (FTMT_F2P_TRIGACK_2),
    .FTMT_F2P_TRIG_3          (FTMT_F2P_TRIG_3),
    .FTMT_F2P_TRIGACK_3       (FTMT_F2P_TRIGACK_3),
    .FTMT_F2P_DEBUG           (FTMT_F2P_DEBUG),
    .FTMT_P2F_TRIGACK_0       (FTMT_P2F_TRIGACK_0),
    .FTMT_P2F_TRIG_0          (FTMT_P2F_TRIG_0),
    .FTMT_P2F_TRIGACK_1       (FTMT_P2F_TRIGACK_1),
    .FTMT_P2F_TRIG_1          (FTMT_P2F_TRIG_1),
    .FTMT_P2F_TRIGACK_2       (FTMT_P2F_TRIGACK_2),
    .FTMT_P2F_TRIG_2          (FTMT_P2F_TRIG_2),
    .FTMT_P2F_TRIGACK_3       (FTMT_P2F_TRIGACK_3),
    .FTMT_P2F_TRIG_3          (FTMT_P2F_TRIG_3),
    .FTMT_P2F_DEBUG           (FTMT_P2F_DEBUG),
  `endif

  `ifdef USE_WATCHDOG
    .WDT_CLK_IN               (WDT_CLK_IN),
    .WDT_RST_OUT              (WDT_RST_OUT),
  `endif
  `ifdef USE_USB0
    .USB0_PORT_INDCTL         (USB0_PORT_INDCTL),
    .USB0_VBUS_PWRSELECT      (USB0_VBUS_PWRSELECT),
    .USB0_VBUS_PWRFAULT       (USB0_VBUS_PWRFAULT),
  `endif
  `ifdef USE_USB1
    .USB1_PORT_INDCTL         (USB1_PORT_INDCTL),
    .USB1_VBUS_PWRSELECT      (USB1_VBUS_PWRSELECT),
    .USB1_VBUS_PWRFAULT       (USB1_VBUS_PWRFAULT),
  `endif
  `ifdef USE_INTERRUPTS
    .IRQ_P2F_DMAC_ABORT       (IRQ_P2F_DMAC_ABORT),
    .IRQ_P2F_DMAC0            (IRQ_P2F_DMAC0),
    .IRQ_P2F_DMAC1            (IRQ_P2F_DMAC1),
    .IRQ_P2F_DMAC2            (IRQ_P2F_DMAC2),
    .IRQ_P2F_DMAC3            (IRQ_P2F_DMAC3),
    .IRQ_P2F_DMAC4            (IRQ_P2F_DMAC4),
    .IRQ_P2F_DMAC5            (IRQ_P2F_DMAC5),
    .IRQ_P2F_DMAC6            (IRQ_P2F_DMAC6),
    .IRQ_P2F_DMAC7            (IRQ_P2F_DMAC7),
    .IRQ_P2F_SMC              (IRQ_P2F_SMC),
    .IRQ_P2F_QSPI             (IRQ_P2F_QSPI),
    .IRQ_P2F_CTI              (IRQ_P2F_CTI),
    .IRQ_P2F_GPIO             (IRQ_P2F_GPIO),
    .IRQ_P2F_USB0             (IRQ_P2F_USB0),
    .IRQ_P2F_ENET0            (IRQ_P2F_ENET0),
    .IRQ_P2F_ENET_WAKE0       (IRQ_P2F_ENET_WAKE0),
    .IRQ_P2F_SDIO0            (IRQ_P2F_SDIO0),
    .IRQ_P2F_I2C0             (IRQ_P2F_I2C0),
    .IRQ_P2F_SPI0             (IRQ_P2F_SPI0),
    .IRQ_P2F_UART0            (IRQ_P2F_UART0),
    .IRQ_P2F_CAN0             (IRQ_P2F_CAN0),
    .IRQ_P2F_USB1             (IRQ_P2F_USB1),
    .IRQ_P2F_ENET1            (IRQ_P2F_ENET1),
    .IRQ_P2F_ENET_WAKE1       (IRQ_P2F_ENET_WAKE1),
    .IRQ_P2F_SDIO1            (IRQ_P2F_SDIO1),
    .IRQ_P2F_I2C1             (IRQ_P2F_I2C1),
    .IRQ_P2F_SPI1             (IRQ_P2F_SPI1),
    .IRQ_P2F_UART1            (IRQ_P2F_UART1),
    .IRQ_P2F_CAN1             (IRQ_P2F_CAN1),
    .Core0_nFIQ               (Core0_nFIQ),
    .Core0_nIRQ               (Core0_nIRQ),
    .Core1_nFIQ               (Core1_nFIQ),
    .Core1_nIRQ               (Core1_nIRQ),
    .IRQ_F2P                  (IRQ_F2P),
    .SRAM_INTIN               (SRAM_INTIN),
  `endif
  `ifdef USE_PS_EVENTS
    .EVENT_EVENTO             (EVENT_EVENTO),
    .EVENT_EVENTI             (EVENT_EVENTI),   
    .EVENT_STANDBYWFE         (EVENT_STANDBYWFE),
    .EVENT_STANDBYWFI         (EVENT_STANDBYWFI),
  `endif
  `ifdef USE_FPGA_IDLE
    .FPGA_IDLE                (FPGA_IDLE),
  `endif    
  `ifdef USE_FCLK0
    .FCLK0_CLK                (FCLK0_CLK),
    .FCLK0_RESET              (FCLK0_RESET),
  `endif
  `ifdef USE_FCLK1
    .FCLK1_CLK                (FCLK1_CLK),
    .FCLK1_RESET              (FCLK1_RESET),
  `endif
  `ifdef USE_FCLK2
    .FCLK2_CLK                (FCLK2_CLK),
    .FCLK2_RESET              (FCLK2_RESET),
  `endif
  `ifdef USE_FCLK3
    .FCLK3_CLK                (FCLK3_CLK),
    .FCLK3_RESET              (FCLK3_RESET),
  `endif
  `ifdef PS_MASTER_AXI_GP0
    .M_AXI_GP0_ACLK           (M_AXI_GP0_clk),
    .M_AXI_GP0_ARESET         (M_AXI_GP0_reset),

    .M_AXI_GP0_ARVALID        (M_AXI_GP0_ar_valid),
    .M_AXI_GP0_AWVALID        (M_AXI_GP0_aw_valid),
    .M_AXI_GP0_BREADY         (M_AXI_GP0_b_ready),
    .M_AXI_GP0_RREADY         (M_AXI_GP0_r_ready),
    .M_AXI_GP0_ARREADY        (M_AXI_GP0_ar_ready),
    .M_AXI_GP0_AWREADY        (M_AXI_GP0_aw_ready),
    .M_AXI_GP0_BVALID         (M_AXI_GP0_b_valid),
    .M_AXI_GP0_RVALID         (M_AXI_GP0_r_valid),
    .M_AXI_GP0_WREADY         (M_AXI_GP0_w_ready),
    .M_AXI_GP0_WVALID         (M_AXI_GP0_w_valid),

    .M_AXI_GP0_WLAST          (M_AXI_GP0_w_payload_last),
    .M_AXI_GP0_ARID           (M_AXI_GP0_ar_payload_id),
    .M_AXI_GP0_AWID           (M_AXI_GP0_aw_payload_id),
    .M_AXI_GP0_WID            (M_AXI_GP0_w_payload_id),
    .M_AXI_GP0_ARBURST        (M_AXI_GP0_ar_payload_burst),
    .M_AXI_GP0_ARLOCK         (M_AXI_GP0_ar_payload_lock_adaptor),
    .M_AXI_GP0_ARSIZE         (M_AXI_GP0_ar_payload_size_adaptor),
    .M_AXI_GP0_AWBURST        (M_AXI_GP0_aw_payload_burst), 
    .M_AXI_GP0_AWLOCK         (M_AXI_GP0_aw_payload_lock_adaptor),
    .M_AXI_GP0_AWSIZE         (M_AXI_GP0_aw_payload_size_adaptor),
    .M_AXI_GP0_ARPROT         (M_AXI_GP0_ar_payload_prot),
    .M_AXI_GP0_AWPROT         (M_AXI_GP0_aw_payload_prot),
    .M_AXI_GP0_ARADDR         (M_AXI_GP0_ar_payload_addr),
    .M_AXI_GP0_AWADDR         (M_AXI_GP0_aw_payload_addr),
    .M_AXI_GP0_WDATA          (M_AXI_GP0_w_payload_data),
    .M_AXI_GP0_ARCACHE        (M_AXI_GP0_ar_payload_cache),
    .M_AXI_GP0_ARLEN          (M_AXI_GP0_ar_payload_len_adaptor),
    .M_AXI_GP0_ARQOS          (M_AXI_GP0_ar_payload_qos),
    .M_AXI_GP0_AWCACHE        (M_AXI_GP0_aw_payload_cache),
    .M_AXI_GP0_AWLEN          (M_AXI_GP0_aw_payload_len_adaptor),
    .M_AXI_GP0_AWQOS          (M_AXI_GP0_aw_payload_qos),
    .M_AXI_GP0_WSTRB          (M_AXI_GP0_w_payload_strb),
    .M_AXI_GP0_RLAST          (M_AXI_GP0_r_payload_last),
    .M_AXI_GP0_BID            (M_AXI_GP0_b_payload_id),
    .M_AXI_GP0_RID            (M_AXI_GP0_r_payload_id),
    .M_AXI_GP0_BRESP          (M_AXI_GP0_b_payload_resp),
    .M_AXI_GP0_RRESP          (M_AXI_GP0_r_payload_resp),
    .M_AXI_GP0_RDATA          (M_AXI_GP0_r_payload_data),  
  `endif
  `ifdef PS_MASTER_AXI_GP1
    .M_AXI_GP1_ACLK           (M_AXI_GP1_ACLK),
    .M_AXI_GP1_ARESET         (M_AXI_GP1_ARESET),
    .M_AXI_GP1_ARVALID        (M_AXI_GP1_ARVALID),
    .M_AXI_GP1_AWVALID        (M_AXI_GP1_AWVALID),
    .M_AXI_GP1_BREADY         (M_AXI_GP1_BREADY),
    .M_AXI_GP1_RREADY         (M_AXI_GP1_RREADY),
    .M_AXI_GP1_WLAST          (M_AXI_GP1_WLAST),
    .M_AXI_GP1_WVALID         (M_AXI_GP1_WVALID),
    .M_AXI_GP1_ARID           (M_AXI_GP1_ARID),
    .M_AXI_GP1_AWID           (M_AXI_GP1_AWID),
    .M_AXI_GP1_WID            (M_AXI_GP1_WID),
    .M_AXI_GP1_ARBURST        (M_AXI_GP1_ARBURST),
    .M_AXI_GP1_ARLOCK         (M_AXI_GP1_ARLOCK),
    .M_AXI_GP1_ARSIZE         (M_AXI_GP1_ARSIZE),
    .M_AXI_GP1_AWBURST        (M_AXI_GP1_AWBURST),
    .M_AXI_GP1_AWLOCK         (M_AXI_GP1_AWLOCK),
    .M_AXI_GP1_AWSIZE         (M_AXI_GP1_AWSIZE),
    .M_AXI_GP1_ARPROT         (M_AXI_GP1_ARPROT),
    .M_AXI_GP1_AWPROT         (M_AXI_GP1_AWPROT),
    .M_AXI_GP1_ARADDR         (M_AXI_GP1_ARADDR),
    .M_AXI_GP1_AWADDR         (M_AXI_GP1_AWADDR),
    .M_AXI_GP1_WDATA          (M_AXI_GP1_WDATA),
    .M_AXI_GP1_ARCACHE        (M_AXI_GP1_ARCACHE),
    .M_AXI_GP1_ARLEN          (M_AXI_GP1_ARLEN),
    .M_AXI_GP1_ARQOS          (M_AXI_GP1_ARQOS),
    .M_AXI_GP1_AWCACHE        (M_AXI_GP1_AWCACHE),
    .M_AXI_GP1_AWLEN          (M_AXI_GP1_AWLEN),
    .M_AXI_GP1_AWQOS          (M_AXI_GP1_AWQOS),
    .M_AXI_GP1_WSTRB          (M_AXI_GP1_WSTRB),
    .M_AXI_GP1_ARREADY        (M_AXI_GP1_ARREADY),
    .M_AXI_GP1_AWREADY        (M_AXI_GP1_AWREADY),
    .M_AXI_GP1_BVALID         (M_AXI_GP1_BVALID),
    .M_AXI_GP1_RLAST          (M_AXI_GP1_RLAST),
    .M_AXI_GP1_RVALID         (M_AXI_GP1_RVALID),
    .M_AXI_GP1_WREADY         (M_AXI_GP1_WREADY),  
    .M_AXI_GP1_BID            (M_AXI_GP1_BID),
    .M_AXI_GP1_RID            (M_AXI_GP1_RID),
    .M_AXI_GP1_BRESP          (M_AXI_GP1_BRESP),
    .M_AXI_GP1_RRESP          (M_AXI_GP1_RRESP),
    .M_AXI_GP1_RDATA          (M_AXI_GP1_RDATA),
  `endif
  `ifdef PS_SLAVE_AXI_GP0
    .S_AXI_GP0_ACLK           (S_AXI_GP0_ACLK),
    .S_AXI_GP0_ARESET         (S_AXI_GP0_ARESET),
    .S_AXI_GP0_ARREADY        (S_AXI_GP0_ARREADY),
    .S_AXI_GP0_AWREADY        (S_AXI_GP0_AWREADY),
    .S_AXI_GP0_BVALID         (S_AXI_GP0_BVALID),
    .S_AXI_GP0_RLAST          (S_AXI_GP0_RLAST),
    .S_AXI_GP0_RVALID         (S_AXI_GP0_RVALID),
    .S_AXI_GP0_WREADY         (S_AXI_GP0_WREADY),  
    .S_AXI_GP0_BRESP          (S_AXI_GP0_BRESP),
    .S_AXI_GP0_RRESP          (S_AXI_GP0_RRESP),
    .S_AXI_GP0_RDATA          (S_AXI_GP0_RDATA),
    .S_AXI_GP0_BID            (S_AXI_GP0_BID),
    .S_AXI_GP0_RID            (S_AXI_GP0_RID),
    .S_AXI_GP0_ARVALID        (S_AXI_GP0_ARVALID),
    .S_AXI_GP0_AWVALID        (S_AXI_GP0_AWVALID),
    .S_AXI_GP0_BREADY         (S_AXI_GP0_BREADY),
    .S_AXI_GP0_RREADY         (S_AXI_GP0_RREADY),
    .S_AXI_GP0_WLAST          (S_AXI_GP0_WLAST),
    .S_AXI_GP0_WVALID         (S_AXI_GP0_WVALID),
    .S_AXI_GP0_ARBURST        (S_AXI_GP0_ARBURST),
    .S_AXI_GP0_ARLOCK         (S_AXI_GP0_ARLOCK),
    .S_AXI_GP0_ARSIZE         (S_AXI_GP0_ARSIZE),
    .S_AXI_GP0_AWBURST        (S_AXI_GP0_AWBURST),
    .S_AXI_GP0_AWLOCK         (S_AXI_GP0_AWLOCK),
    .S_AXI_GP0_AWSIZE         (S_AXI_GP0_AWSIZE),
    .S_AXI_GP0_ARPROT         (S_AXI_GP0_ARPROT),
    .S_AXI_GP0_AWPROT         (S_AXI_GP0_AWPROT),
    .S_AXI_GP0_ARADDR         (S_AXI_GP0_ARADDR),
    .S_AXI_GP0_AWADDR         (S_AXI_GP0_AWADDR),
    .S_AXI_GP0_WDATA          (S_AXI_GP0_WDATA),
    .S_AXI_GP0_ARCACHE        (S_AXI_GP0_ARCACHE),
    .S_AXI_GP0_ARLEN          (S_AXI_GP0_ARLEN),
    .S_AXI_GP0_ARQOS          (S_AXI_GP0_ARQOS),
    .S_AXI_GP0_AWCACHE        (S_AXI_GP0_AWCACHE),
    .S_AXI_GP0_AWLEN          (S_AXI_GP0_AWLEN),
    .S_AXI_GP0_AWQOS          (S_AXI_GP0_AWQOS),
    .S_AXI_GP0_WSTRB          (S_AXI_GP0_WSTRB),
    .S_AXI_GP0_ARID           (S_AXI_GP0_ARID),
    .S_AXI_GP0_AWID           (S_AXI_GP0_AWID),
    .S_AXI_GP0_WID            (S_AXI_GP0_WID), 
  `endif
  `ifdef PS_SLAVE_AXI_GP1
    .S_AXI_GP1_ACLK           (S_AXI_GP1_ACLK),
    .S_AXI_GP1_ARESET         (S_AXI_GP1_ARESET),
    .S_AXI_GP1_ARREADY        (S_AXI_GP1_ARREADY),
    .S_AXI_GP1_AWREADY        (S_AXI_GP1_AWREADY),
    .S_AXI_GP1_BVALID         (S_AXI_GP1_BVALID),
    .S_AXI_GP1_RLAST          (S_AXI_GP1_RLAST),
    .S_AXI_GP1_RVALID         (S_AXI_GP1_RVALID),
    .S_AXI_GP1_WREADY         (S_AXI_GP1_WREADY),  
    .S_AXI_GP1_BRESP          (S_AXI_GP1_BRESP),
    .S_AXI_GP1_RRESP          (S_AXI_GP1_RRESP),
    .S_AXI_GP1_RDATA          (S_AXI_GP1_RDATA),
    .S_AXI_GP1_BID            (S_AXI_GP1_BID),
    .S_AXI_GP1_RID            (S_AXI_GP1_RID),
    .S_AXI_GP1_ARVALID        (S_AXI_GP1_ARVALID),
    .S_AXI_GP1_AWVALID        (S_AXI_GP1_AWVALID),
    .S_AXI_GP1_BREADY         (S_AXI_GP1_BREADY),
    .S_AXI_GP1_RREADY         (S_AXI_GP1_RREADY),
    .S_AXI_GP1_WLAST          (S_AXI_GP1_WLAST),
    .S_AXI_GP1_WVALID         (S_AXI_GP1_WVALID),
    .S_AXI_GP1_ARBURST        (S_AXI_GP1_ARBURST),
    .S_AXI_GP1_ARLOCK         (S_AXI_GP1_ARLOCK),
    .S_AXI_GP1_ARSIZE         (S_AXI_GP1_ARSIZE),
    .S_AXI_GP1_AWBURST        (S_AXI_GP1_AWBURST),
    .S_AXI_GP1_AWLOCK         (S_AXI_GP1_AWLOCK),
    .S_AXI_GP1_AWSIZE         (S_AXI_GP1_AWSIZE),
    .S_AXI_GP1_ARPROT         (S_AXI_GP1_ARPROT),
    .S_AXI_GP1_AWPROT         (S_AXI_GP1_AWPROT),
    .S_AXI_GP1_ARADDR         (S_AXI_GP1_ARADDR),
    .S_AXI_GP1_AWADDR         (S_AXI_GP1_AWADDR),
    .S_AXI_GP1_WDATA          (S_AXI_GP1_WDATA),
    .S_AXI_GP1_ARCACHE        (S_AXI_GP1_ARCACHE),
    .S_AXI_GP1_ARLEN          (S_AXI_GP1_ARLEN),
    .S_AXI_GP1_ARQOS          (S_AXI_GP1_ARQOS),
    .S_AXI_GP1_AWCACHE        (S_AXI_GP1_AWCACHE),
    .S_AXI_GP1_AWLEN          (S_AXI_GP1_AWLEN),
    .S_AXI_GP1_AWQOS          (S_AXI_GP1_AWQOS),
    .S_AXI_GP1_WSTRB          (S_AXI_GP1_WSTRB),
    .S_AXI_GP1_ARID           (S_AXI_GP1_ARID),
    .S_AXI_GP1_AWID           (S_AXI_GP1_AWID),
    .S_AXI_GP1_WID            (S_AXI_GP1_WID), 
  `endif
  `ifdef PS_SLAVE_AXI_ACP
    .S_AXI_ACP_ACLK           (S_AXI_ACP_ACLK),
    .S_AXI_ACP_ARESET         (S_AXI_ACP_ARESET),
    .S_AXI_ACP_ARREADY        (S_AXI_ACP_ARREADY),
    .S_AXI_ACP_AWREADY        (S_AXI_ACP_AWREADY),
    .S_AXI_ACP_BVALID         (S_AXI_ACP_BVALID),
    .S_AXI_ACP_RLAST          (S_AXI_ACP_RLAST),
    .S_AXI_ACP_RVALID         (S_AXI_ACP_RVALID),
    .S_AXI_ACP_WREADY         (S_AXI_ACP_WREADY),  
    .S_AXI_ACP_BRESP          (S_AXI_ACP_BRESP),
    .S_AXI_ACP_RRESP          (S_AXI_ACP_RRESP),
    .S_AXI_ACP_BID            (S_AXI_ACP_BID),
    .S_AXI_ACP_RID            (S_AXI_ACP_RID),
    .S_AXI_ACP_RDATA          (S_AXI_ACP_RDATA),
    .S_AXI_ACP_ARVALID        (S_AXI_ACP_ARVALID),
    .S_AXI_ACP_AWVALID        (S_AXI_ACP_AWVALID),
    .S_AXI_ACP_BREADY         (S_AXI_ACP_BREADY),
    .S_AXI_ACP_RREADY         (S_AXI_ACP_RREADY),
    .S_AXI_ACP_WLAST          (S_AXI_ACP_WLAST),
    .S_AXI_ACP_WVALID         (S_AXI_ACP_WVALID),
    .S_AXI_ACP_ARID           (S_AXI_ACP_ARID),
    .S_AXI_ACP_ARPROT         (S_AXI_ACP_ARPROT),
    .S_AXI_ACP_AWID           (S_AXI_ACP_AWID),
    .S_AXI_ACP_AWPROT         (S_AXI_ACP_AWPROT),
    .S_AXI_ACP_WID            (S_AXI_ACP_WID),
    .S_AXI_ACP_ARADDR         (S_AXI_ACP_ARADDR),
    .S_AXI_ACP_AWADDR         (S_AXI_ACP_AWADDR),
    .S_AXI_ACP_ARCACHE        (S_AXI_ACP_ARCACHE),
    .S_AXI_ACP_ARLEN          (S_AXI_ACP_ARLEN),
    .S_AXI_ACP_ARQOS          (S_AXI_ACP_ARQOS),
    .S_AXI_ACP_AWCACHE        (S_AXI_ACP_AWCACHE),
    .S_AXI_ACP_AWLEN          (S_AXI_ACP_AWLEN),
    .S_AXI_ACP_AWQOS          (S_AXI_ACP_AWQOS),
    .S_AXI_ACP_ARBURST        (S_AXI_ACP_ARBURST),
    .S_AXI_ACP_ARLOCK         (S_AXI_ACP_ARLOCK),
    .S_AXI_ACP_ARSIZE         (S_AXI_ACP_ARSIZE),
    .S_AXI_ACP_AWBURST        (S_AXI_ACP_AWBURST),
    .S_AXI_ACP_AWLOCK         (S_AXI_ACP_AWLOCK),
    .S_AXI_ACP_AWSIZE         (S_AXI_ACP_AWSIZE),
    .S_AXI_ACP_ARUSER         (S_AXI_ACP_ARUSER),
    .S_AXI_ACP_AWUSER         (S_AXI_ACP_AWUSER),
    .S_AXI_ACP_WDATA          (S_AXI_ACP_WDATA),
    .S_AXI_ACP_WSTRB          (S_AXI_ACP_WSTRB), 
  `endif
  `ifdef PS_SLAVE_AXI_HP0
    .S_AXI_HP0_ARESET         (S_AXI_HP0_ARESET),
    .S_AXI_HP0_ARREADY        (S_AXI_HP0_ARREADY),
    .S_AXI_HP0_AWREADY        (S_AXI_HP0_AWREADY),
    .S_AXI_HP0_BVALID         (S_AXI_HP0_BVALID),
    .S_AXI_HP0_RLAST          (S_AXI_HP0_RLAST),
    .S_AXI_HP0_RVALID         (S_AXI_HP0_RVALID),
    .S_AXI_HP0_WREADY         (S_AXI_HP0_WREADY),  
    .S_AXI_HP0_BRESP          (S_AXI_HP0_BRESP),
    .S_AXI_HP0_RRESP          (S_AXI_HP0_RRESP),
    .S_AXI_HP0_BID            (S_AXI_HP0_BID),
    .S_AXI_HP0_RID            (S_AXI_HP0_RID),
    .S_AXI_HP0_RDATA          (S_AXI_HP0_RDATA),
    .S_AXI_HP0_RCOUNT         (S_AXI_HP0_RCOUNT),
    .S_AXI_HP0_WCOUNT         (S_AXI_HP0_WCOUNT),
    .S_AXI_HP0_RACOUNT        (S_AXI_HP0_RACOUNT),
    .S_AXI_HP0_WACOUNT        (S_AXI_HP0_WACOUNT),
    .S_AXI_HP0_ACLK           (S_AXI_HP0_ACLK),
    .S_AXI_HP0_ARVALID        (S_AXI_HP0_ARVALID),
    .S_AXI_HP0_AWVALID        (S_AXI_HP0_AWVALID),
    .S_AXI_HP0_BREADY         (S_AXI_HP0_BREADY),
    .S_AXI_HP0_RDISSUECAP1_EN (S_AXI_HP0_RDISSUECAP1_EN),
    .S_AXI_HP0_RREADY         (S_AXI_HP0_RREADY),
    .S_AXI_HP0_WLAST          (S_AXI_HP0_WLAST),
    .S_AXI_HP0_WRISSUECAP1_EN (S_AXI_HP0_WRISSUECAP1_EN),
    .S_AXI_HP0_WVALID         (S_AXI_HP0_WVALID),
    .S_AXI_HP0_ARBURST        (S_AXI_HP0_ARBURST),
    .S_AXI_HP0_ARLOCK         (S_AXI_HP0_ARLOCK),
    .S_AXI_HP0_ARSIZE         (S_AXI_HP0_ARSIZE),
    .S_AXI_HP0_AWBURST        (S_AXI_HP0_AWBURST),
    .S_AXI_HP0_AWLOCK         (S_AXI_HP0_AWLOCK),
    .S_AXI_HP0_AWSIZE         (S_AXI_HP0_AWSIZE),
    .S_AXI_HP0_ARPROT         (S_AXI_HP0_ARPROT),
    .S_AXI_HP0_AWPROT         (S_AXI_HP0_AWPROT),
    .S_AXI_HP0_ARADDR         (S_AXI_HP0_ARADDR),
    .S_AXI_HP0_AWADDR         (S_AXI_HP0_AWADDR),
    .S_AXI_HP0_ARCACHE        (S_AXI_HP0_ARCACHE),
    .S_AXI_HP0_ARLEN          (S_AXI_HP0_ARLEN),
    .S_AXI_HP0_ARQOS          (S_AXI_HP0_ARQOS),
    .S_AXI_HP0_AWCACHE        (S_AXI_HP0_AWCACHE),
    .S_AXI_HP0_AWLEN          (S_AXI_HP0_AWLEN),
    .S_AXI_HP0_AWQOS          (S_AXI_HP0_AWQOS),
    .S_AXI_HP0_ARID           (S_AXI_HP0_ARID),
    .S_AXI_HP0_AWID           (S_AXI_HP0_AWID),
    .S_AXI_HP0_WID            (S_AXI_HP0_WID),
    .S_AXI_HP0_WDATA          (S_AXI_HP0_WDATA),
    .S_AXI_HP0_WSTRB          (S_AXI_HP0_WSTRB),
  `endif
  `ifdef PS_SLAVE_AXI_HP1
    .S_AXI_HP1_ARESET         (S_AXI_HP1_ARESET),
    .S_AXI_HP1_ARREADY        (S_AXI_HP1_ARREADY),
    .S_AXI_HP1_AWREADY        (S_AXI_HP1_AWREADY),
    .S_AXI_HP1_BVALID         (S_AXI_HP1_BVALID),
    .S_AXI_HP1_RLAST          (S_AXI_HP1_RLAST),
    .S_AXI_HP1_RVALID         (S_AXI_HP1_RVALID),
    .S_AXI_HP1_WREADY         (S_AXI_HP1_WREADY),  
    .S_AXI_HP1_BRESP          (S_AXI_HP1_BRESP),
    .S_AXI_HP1_RRESP          (S_AXI_HP1_RRESP),
    .S_AXI_HP1_BID            (S_AXI_HP1_BID),
    .S_AXI_HP1_RID            (S_AXI_HP1_RID),
    .S_AXI_HP1_RDATA          (S_AXI_HP1_RDATA),
    .S_AXI_HP1_RCOUNT         (S_AXI_HP1_RCOUNT),
    .S_AXI_HP1_WCOUNT         (S_AXI_HP1_WCOUNT),
    .S_AXI_HP1_RACOUNT        (S_AXI_HP1_RACOUNT),
    .S_AXI_HP1_WACOUNT        (S_AXI_HP1_WACOUNT),
    .S_AXI_HP1_ACLK           (S_AXI_HP1_ACLK),
    .S_AXI_HP1_ARVALID        (S_AXI_HP1_ARVALID),
    .S_AXI_HP1_AWVALID        (S_AXI_HP1_AWVALID),
    .S_AXI_HP1_BREADY         (S_AXI_HP1_BREADY),
    .S_AXI_HP1_RDISSUECAP1_EN (S_AXI_HP1_RDISSUECAP1_EN),
    .S_AXI_HP1_RREADY         (S_AXI_HP1_RREADY),
    .S_AXI_HP1_WLAST          (S_AXI_HP1_WLAST),
    .S_AXI_HP1_WRISSUECAP1_EN (S_AXI_HP1_WRISSUECAP1_EN),
    .S_AXI_HP1_WVALID         (S_AXI_HP1_WVALID),
    .S_AXI_HP1_ARBURST        (S_AXI_HP1_ARBURST),
    .S_AXI_HP1_ARLOCK         (S_AXI_HP1_ARLOCK),
    .S_AXI_HP1_ARSIZE         (S_AXI_HP1_ARSIZE),
    .S_AXI_HP1_AWBURST        (S_AXI_HP1_AWBURST),
    .S_AXI_HP1_AWLOCK         (S_AXI_HP1_AWLOCK),
    .S_AXI_HP1_AWSIZE         (S_AXI_HP1_AWSIZE),
    .S_AXI_HP1_ARPROT         (S_AXI_HP1_ARPROT),
    .S_AXI_HP1_AWPROT         (S_AXI_HP1_AWPROT),
    .S_AXI_HP1_ARADDR         (S_AXI_HP1_ARADDR),
    .S_AXI_HP1_AWADDR         (S_AXI_HP1_AWADDR),
    .S_AXI_HP1_ARCACHE        (S_AXI_HP1_ARCACHE),
    .S_AXI_HP1_ARLEN          (S_AXI_HP1_ARLEN),
    .S_AXI_HP1_ARQOS          (S_AXI_HP1_ARQOS),
    .S_AXI_HP1_AWCACHE        (S_AXI_HP1_AWCACHE),
    .S_AXI_HP1_AWLEN          (S_AXI_HP1_AWLEN),
    .S_AXI_HP1_AWQOS          (S_AXI_HP1_AWQOS),
    .S_AXI_HP1_ARID           (S_AXI_HP1_ARID),
    .S_AXI_HP1_AWID           (S_AXI_HP1_AWID),
    .S_AXI_HP1_WID            (S_AXI_HP1_WID),
    .S_AXI_HP1_WDATA          (S_AXI_HP1_WDATA),
    .S_AXI_HP1_WSTRB          (S_AXI_HP1_WSTRB),
  `endif
  `ifdef PS_SLAVE_AXI_HP2
    .S_AXI_HP2_ARESET         (S_AXI_HP2_ARESET),
    .S_AXI_HP2_ARREADY        (S_AXI_HP2_ARREADY),
    .S_AXI_HP2_AWREADY        (S_AXI_HP2_AWREADY),
    .S_AXI_HP2_BVALID         (S_AXI_HP2_BVALID),
    .S_AXI_HP2_RLAST          (S_AXI_HP2_RLAST),
    .S_AXI_HP2_RVALID         (S_AXI_HP2_RVALID),
    .S_AXI_HP2_WREADY         (S_AXI_HP2_WREADY),  
    .S_AXI_HP2_BRESP          (S_AXI_HP2_BRESP),
    .S_AXI_HP2_RRESP          (S_AXI_HP2_RRESP),
    .S_AXI_HP2_BID            (S_AXI_HP2_BID),
    .S_AXI_HP2_RID            (S_AXI_HP2_RID),
    .S_AXI_HP2_RDATA          (S_AXI_HP2_RDATA),
    .S_AXI_HP2_RCOUNT         (S_AXI_HP2_RCOUNT),
    .S_AXI_HP2_WCOUNT         (S_AXI_HP2_WCOUNT),
    .S_AXI_HP2_RACOUNT        (S_AXI_HP2_RACOUNT),
    .S_AXI_HP2_WACOUNT        (S_AXI_HP2_WACOUNT),
    .S_AXI_HP2_ACLK           (S_AXI_HP2_ACLK),
    .S_AXI_HP2_ARVALID        (S_AXI_HP2_ARVALID),
    .S_AXI_HP2_AWVALID        (S_AXI_HP2_AWVALID),
    .S_AXI_HP2_BREADY         (S_AXI_HP2_BREADY),
    .S_AXI_HP2_RDISSUECAP1_EN (S_AXI_HP2_RDISSUECAP1_EN),
    .S_AXI_HP2_RREADY         (S_AXI_HP2_RREADY),
    .S_AXI_HP2_WLAST          (S_AXI_HP2_WLAST),
    .S_AXI_HP2_WRISSUECAP1_EN (S_AXI_HP2_WRISSUECAP1_EN),
    .S_AXI_HP2_WVALID         (S_AXI_HP2_WVALID),
    .S_AXI_HP2_ARBURST        (S_AXI_HP2_ARBURST),
    .S_AXI_HP2_ARLOCK         (S_AXI_HP2_ARLOCK),
    .S_AXI_HP2_ARSIZE         (S_AXI_HP2_ARSIZE),
    .S_AXI_HP2_AWBURST        (S_AXI_HP2_AWBURST),
    .S_AXI_HP2_AWLOCK         (S_AXI_HP2_AWLOCK),
    .S_AXI_HP2_AWSIZE         (S_AXI_HP2_AWSIZE),
    .S_AXI_HP2_ARPROT         (S_AXI_HP2_ARPROT),
    .S_AXI_HP2_AWPROT         (S_AXI_HP2_AWPROT),
    .S_AXI_HP2_ARADDR         (S_AXI_HP2_ARADDR),
    .S_AXI_HP2_AWADDR         (S_AXI_HP2_AWADDR),
    .S_AXI_HP2_ARCACHE        (S_AXI_HP2_ARCACHE),
    .S_AXI_HP2_ARLEN          (S_AXI_HP2_ARLEN),
    .S_AXI_HP2_ARQOS          (S_AXI_HP2_ARQOS),
    .S_AXI_HP2_AWCACHE        (S_AXI_HP2_AWCACHE),
    .S_AXI_HP2_AWLEN          (S_AXI_HP2_AWLEN),
    .S_AXI_HP2_AWQOS          (S_AXI_HP2_AWQOS),
    .S_AXI_HP2_ARID           (S_AXI_HP2_ARID),
    .S_AXI_HP2_AWID           (S_AXI_HP2_AWID),
    .S_AXI_HP2_WID            (S_AXI_HP2_WID),
    .S_AXI_HP2_WDATA          (S_AXI_HP2_WDATA),
    .S_AXI_HP2_WSTRB          (S_AXI_HP2_WSTRB),
  `endif
  `ifdef PS_SLAVE_AXI_HP3
    .S_AXI_HP3_ARESET         (S_AXI_HP3_ARESET),
    .S_AXI_HP3_ARREADY        (S_AXI_HP3_ARREADY),
    .S_AXI_HP3_AWREADY        (S_AXI_HP3_AWREADY),
    .S_AXI_HP3_BVALID         (S_AXI_HP3_BVALID),
    .S_AXI_HP3_RLAST          (S_AXI_HP3_RLAST),
    .S_AXI_HP3_RVALID         (S_AXI_HP3_RVALID),
    .S_AXI_HP3_WREADY         (S_AXI_HP3_WREADY),  
    .S_AXI_HP3_BRESP          (S_AXI_HP3_BRESP),
    .S_AXI_HP3_RRESP          (S_AXI_HP3_RRESP),
    .S_AXI_HP3_BID            (S_AXI_HP3_BID),
    .S_AXI_HP3_RID            (S_AXI_HP3_RID),
    .S_AXI_HP3_RDATA          (S_AXI_HP3_RDATA),
    .S_AXI_HP3_RCOUNT         (S_AXI_HP3_RCOUNT),
    .S_AXI_HP3_WCOUNT         (S_AXI_HP3_WCOUNT),
    .S_AXI_HP3_RACOUNT        (S_AXI_HP3_RACOUNT),
    .S_AXI_HP3_WACOUNT        (S_AXI_HP3_WACOUNT),
    .S_AXI_HP3_ACLK           (S_AXI_HP3_ACLK),
    .S_AXI_HP3_ARVALID        (S_AXI_HP3_ARVALID),
    .S_AXI_HP3_AWVALID        (S_AXI_HP3_AWVALID),
    .S_AXI_HP3_BREADY         (S_AXI_HP3_BREADY),
    .S_AXI_HP3_RDISSUECAP1_EN (S_AXI_HP3_RDISSUECAP1_EN),
    .S_AXI_HP3_RREADY         (S_AXI_HP3_RREADY),
    .S_AXI_HP3_WLAST          (S_AXI_HP3_WLAST),
    .S_AXI_HP3_WRISSUECAP1_EN (S_AXI_HP3_WRISSUECAP1_EN),
    .S_AXI_HP3_WVALID         (S_AXI_HP3_WVALID),
    .S_AXI_HP3_ARBURST        (S_AXI_HP3_ARBURST),
    .S_AXI_HP3_ARLOCK         (S_AXI_HP3_ARLOCK),
    .S_AXI_HP3_ARSIZE         (S_AXI_HP3_ARSIZE),
    .S_AXI_HP3_AWBURST        (S_AXI_HP3_AWBURST),
    .S_AXI_HP3_AWLOCK         (S_AXI_HP3_AWLOCK),
    .S_AXI_HP3_AWSIZE         (S_AXI_HP3_AWSIZE),
    .S_AXI_HP3_ARPROT         (S_AXI_HP3_ARPROT),
    .S_AXI_HP3_AWPROT         (S_AXI_HP3_AWPROT),
    .S_AXI_HP3_ARADDR         (S_AXI_HP3_ARADDR),
    .S_AXI_HP3_AWADDR         (S_AXI_HP3_AWADDR),
    .S_AXI_HP3_ARCACHE        (S_AXI_HP3_ARCACHE),
    .S_AXI_HP3_ARLEN          (S_AXI_HP3_ARLEN),
    .S_AXI_HP3_ARQOS          (S_AXI_HP3_ARQOS),
    .S_AXI_HP3_AWCACHE        (S_AXI_HP3_AWCACHE),
    .S_AXI_HP3_AWLEN          (S_AXI_HP3_AWLEN),
    .S_AXI_HP3_AWQOS          (S_AXI_HP3_AWQOS),
    .S_AXI_HP3_ARID           (S_AXI_HP3_ARID),
    .S_AXI_HP3_AWID           (S_AXI_HP3_AWID),
    .S_AXI_HP3_WID            (S_AXI_HP3_WID),
    .S_AXI_HP3_WDATA          (S_AXI_HP3_WDATA),
    .S_AXI_HP3_WSTRB          (S_AXI_HP3_WSTRB),
  `endif
  // DDR
  .DDR_ARB                  (DDR_ARB),
  .DDR_CAS_n                (DDR_CAS_n),
  .DDR_CKE                  (DDR_CKE),
  .DDR_Clk_n                (DDR_Clk_n),
  .DDR_Clk                  (DDR_Clk),
  .DDR_CS_n                 (DDR_CS_n),
  .DDR_DRSTB                (DDR_DRSTB),
  .DDR_ODT                  (DDR_ODT),
  .DDR_RAS_n                (DDR_RAS_n),
  .DDR_WEB                  (DDR_WEB),
  .DDR_BankAddr             (DDR_BankAddr),
  .DDR_Addr                 (DDR_Addr),
  .DDR_VRN                  (DDR_VRN),
  .DDR_VRP                  (DDR_VRP),
  .DDR_DM                   (DDR_DM),
  .DDR_DQ                   (DDR_DQ),
  .DDR_DQS_n                (DDR_DQS_n),
  .DDR_DQS                  (DDR_DQS),
  // PS Clock and Reset wires
  .PS_CLK                   (PS_CLK),         
  .PS_SYSTEM_RESET          (PS_SYSTEM_RESET),
  .PS_POWER_ON_RESET        (PS_POWER_ON_RESET)

  );
endmodule
