
module ps7_port_rename( 
  //CAN wires
  output wire CAN0_PHY_TX,
  input wire CAN0_PHY_RX,
  output wire CAN1_PHY_TX,  
  input wire  CAN1_PHY_RX,
  
  //Ethernet wires
  output wire ENET0_GMII_TX_EN,
  output wire ENET0_GMII_TX_ER,
  output wire ENET0_MDIO_MDC,
  output wire ENET0_MDIO_O,
  output wire ENET0_MDIO_T_n,
  output wire ENET0_PTP_DELAY_REQ_RX,
  output wire ENET0_PTP_DELAY_REQ_TX,
  output wire ENET0_PTP_PDELAY_REQ_RX,
  output wire ENET0_PTP_PDELAY_REQ_TX,
  output wire ENET0_PTP_PDELAY_RESP_RX,
  output wire ENET0_PTP_PDELAY_RESP_TX,
  output wire ENET0_PTP_SYNC_FRAME_RX,
  output wire ENET0_PTP_SYNC_FRAME_TX,
  output wire ENET0_SOF_RX,
  output wire ENET0_SOF_TX,
  output wire [7:0] ENET0_GMII_TXD,  
  input wire ENET0_GMII_COL,
  input wire ENET0_GMII_CRS,
  input wire ENET0_GMII_RX_CLK,
  input wire ENET0_GMII_RX_DV,
  input wire ENET0_GMII_RX_ER,
  input wire ENET0_GMII_TX_CLK,
  input wire ENET0_MDIO_I,
  input wire ENET0_EXT_INTIN,
  input wire [7:0] ENET0_GMII_RXD,  

  output wire ENET1_GMII_TX_EN,
  output wire ENET1_GMII_TX_ER,
  output wire ENET1_MDIO_MDC,
  output wire ENET1_MDIO_O,
  output wire ENET1_MDIO_T_n,
  output wire ENET1_PTP_DELAY_REQ_RX,
  output wire ENET1_PTP_DELAY_REQ_TX,
  output wire ENET1_PTP_PDELAY_REQ_RX,
  output wire ENET1_PTP_PDELAY_REQ_TX,
  output wire ENET1_PTP_PDELAY_RESP_RX,
  output wire ENET1_PTP_PDELAY_RESP_TX,
  output wire ENET1_PTP_SYNC_FRAME_RX,
  output wire ENET1_PTP_SYNC_FRAME_TX,
  output wire ENET1_SOF_RX,
  output wire ENET1_SOF_TX,
  output wire [7:0] ENET1_GMII_TXD,
  input wire ENET1_GMII_COL,
  input wire ENET1_GMII_CRS,
  input wire ENET1_GMII_RX_CLK,
  input wire ENET1_GMII_RX_DV,
  input wire ENET1_GMII_RX_ER,
  input wire ENET1_GMII_TX_CLK,
  input wire ENET1_MDIO_I,
  input wire ENET1_EXT_INTIN,  
  input wire [7:0] ENET1_GMII_RXD,

  // 4 DMA ports
  input wire DMA0_ACLK,
  output wire DMA0_RESET_n,  
  output wire [1:0] DMA0_DATYPE,  
  input wire [1:0] DMA0_DRTYPE,
  output wire DMA0_DAVALID,
  output wire DMA0_DRREADY,
  input wire DMA0_DAREADY,
  input wire DMA0_DRLAST,
  input wire DMA0_DRVALID,

  input wire DMA1_ACLK,
  output wire DMA1_RESET_n,  
  output wire [1:0] DMA1_DATYPE,  
  input wire [1:0] DMA1_DRTYPE,
  output wire DMA1_DAVALID,
  output wire DMA1_DRREADY,
  input wire DMA1_DAREADY,
  input wire DMA1_DRLAST,
  input wire DMA1_DRVALID,

  input wire DMA2_ACLK,
  output wire DMA2_RESET_n,  
  output wire [1:0] DMA2_DATYPE,  
  input wire [1:0] DMA2_DRTYPE,
  output wire DMA2_DAVALID,
  output wire DMA2_DRREADY,
  input wire DMA2_DAREADY,
  input wire DMA2_DRLAST,
  input wire DMA2_DRVALID,

  input wire DMA3_ACLK,
  output wire DMA3_RESET_n,  
  output wire [1:0] DMA3_DATYPE,    
  input wire [1:0] DMA3_DRTYPE,
  output wire DMA3_DRREADY,
  input wire DMA3_DAREADY,
  input wire DMA3_DRLAST,
  input wire DMA3_DRVALID,  
  output wire DMA3_DAVALID,

  // tristate GPIO wires + 54 MIO
  input wire [63:0] GPIO_I,
  output wire [63:0] GPIO_O,
  output wire [63:0] GPIO_T_n,
  inout wire [53:0] MIO,  
  
  //I2C wires
  input wire I2C0_SDA_I,
  output wire I2C0_SDA_O,
  output wire I2C0_SDA_T_n,
  input wire I2C0_SCL_I,
  output wire I2C0_SCL_O,
  output wire I2C0_SCL_T_n,
  
  input wire I2C1_SDA_I,
  output wire I2C1_SDA_O,
  output wire I2C1_SDA_T_n,
  input wire I2C1_SCL_I,
  output wire I2C1_SCL_O,
  output wire I2C1_SCL_T_n,
   
  //SDIO wires
  output wire SDIO0_CLK,
  input wire SDIO0_CLK_FB,
  output wire SDIO0_CMD_O,
  input wire SDIO0_CMD_I,
  output wire SDIO0_CMD_T_n,
  input wire [3:0] SDIO0_DATA_I,
  output wire [3:0] SDIO0_DATA_O,
  output wire [3:0] SDIO0_DATA_T_n,
  output wire SDIO0_LED,
  input wire SDIO0_CDN,
  input wire SDIO0_WP,  
  output wire SDIO0_BUSPOW,
  output wire [2:0] SDIO0_BUSVOLT,
  output wire SDIO1_CLK,
  input wire SDIO1_CLK_FB,
  output wire SDIO1_CMD_O,
  input wire SDIO1_CMD_I,
  output wire SDIO1_CMD_T_n,
  input wire [3:0] SDIO1_DATA_I,
  output wire [3:0] SDIO1_DATA_O,
  output wire [3:0] SDIO1_DATA_T_n,
  output wire SDIO1_LED,
  input wire SDIO1_CDN,
  input wire SDIO1_WP,
  output wire SDIO1_BUSPOW,
  output wire [2:0] SDIO1_BUSVOLT,

  // SPI wires
  input wire SPI0_SCLK_I,
  output  wire SPI0_SCLK_O,
  output wire SPI0_SCLK_T_n,
  input wire SPI0_MOSI_I,
  output wire SPI0_MOSI_O,
  output wire SPI0_MOSI_T_n,
  input wire SPI0_MISO_I,
  output wire SPI0_MISO_O,
  output wire SPI0_MISO_T_n,
  input wire SPI0_SS_I,
  output wire SPI0_SS_O,
  output wire SPI0_SS1_O,
  output wire SPI0_SS2_O,
  output wire SPI0_SS_T_n,
  input wire SPI1_SCLK_I,
  output wire SPI1_SCLK_O,
  output wire SPI1_SCLK_T_n,
  input wire SPI1_MOSI_I,
  output wire SPI1_MOSI_O,
  output wire SPI1_MOSI_T_n,
  input wire SPI1_MISO_I,
  output wire SPI1_MISO_O,
  output wire SPI1_MISO_T_n,
  input wire SPI1_SS_I,
  output wire SPI1_SS_O,
  output wire SPI1_SS1_O,
  output wire SPI1_SS2_O,
  output wire SPI1_SS_T_n,

  // UART wires
  output wire UART0_DTRN,
  output wire UART0_RTSN, 
  output wire UART0_TX,
  input wire UART0_CTSN,
  input wire UART0_DCDN,
  input wire UART0_DSRN,
  input wire UART0_RIN,
  input wire UART0_RX,
  output wire UART1_DTRN,
  output wire UART1_RTSN,  
  output wire UART1_TX,
  input wire UART1_CTSN,
  input wire UART1_DCDN,
  input wire UART1_DSRN,
  input wire UART1_RIN,
  input wire UART1_RX,

  //JTAG and trace wires
  input wire PJTAG_TCK,
  input wire PJTAG_TMS,
  input wire PJTAG_TDI,
  output wire PJTAG_TDO_O,
  output wire PJTAG_TDO_T_n,
  output wire TTC0_WAVE0_OUT,
  output wire TTC0_WAVE1_OUT,
  output wire TTC0_WAVE2_OUT,
  input wire TTC0_CLK0_IN,
  input wire TTC0_CLK1_IN,
  input wire TTC0_CLK2_IN,
  output wire TTC1_WAVE0_OUT,
  output wire TTC1_WAVE1_OUT,
  output wire TTC1_WAVE2_OUT,
  input wire TTC1_CLK0_IN,
  input wire TTC1_CLK1_IN,
  input wire TTC1_CLK2_IN,
  input wire TRACE_CLK,
  output wire TRACE_CTL,
  output wire [31:0] TRACE_DATA,
  output wire TRACE_CLK_OUT,
  input wire [31:0] FTMD_TRACEIN_DATA,
  input wire FTMD_TRACEIN_VALID,
  input wire FTMD_TRACEIN_CLK,
  input wire [3:0]  FTMD_TRACEIN_ATID,
  input wire FTMT_F2P_TRIG_0,
  output wire FTMT_F2P_TRIGACK_0,
  input wire FTMT_F2P_TRIG_1,
  output wire FTMT_F2P_TRIGACK_1,
  input wire FTMT_F2P_TRIG_2,
  output wire FTMT_F2P_TRIGACK_2,
  input wire FTMT_F2P_TRIG_3,
  output wire FTMT_F2P_TRIGACK_3,
  input wire [31:0] FTMT_F2P_DEBUG,
  input wire FTMT_P2F_TRIGACK_0,
  output wire FTMT_P2F_TRIG_0,
  input wire FTMT_P2F_TRIGACK_1,
  output wire FTMT_P2F_TRIG_1,
  input wire FTMT_P2F_TRIGACK_2,
  output wire FTMT_P2F_TRIG_2,
  input wire FTMT_P2F_TRIGACK_3,
  output wire FTMT_P2F_TRIG_3,
  output wire [31:0] FTMT_P2F_DEBUG,

  // Watchdog wires
  input wire WDT_CLK_IN,
  output wire WDT_RST_OUT,
 
  // USB wires
  output wire [1:0] USB0_PORT_INDCTL,
  output wire USB0_VBUS_PWRSELECT,
  input wire USB0_VBUS_PWRFAULT,
  output wire [1:0]  USB1_PORT_INDCTL,
  output wire USB1_VBUS_PWRSELECT,
  input wire USB1_VBUS_PWRFAULT,
  
  input wire SRAM_INTIN,

  // events and interrupts
  output wire IRQ_P2F_DMAC_ABORT,
  output wire IRQ_P2F_DMAC0,
  output wire IRQ_P2F_DMAC1,
  output wire IRQ_P2F_DMAC2,
  output wire IRQ_P2F_DMAC3,
  output wire IRQ_P2F_DMAC4,
  output wire IRQ_P2F_DMAC5,
  output wire IRQ_P2F_DMAC6,
  output wire IRQ_P2F_DMAC7,
  output wire IRQ_P2F_SMC,
  output wire IRQ_P2F_QSPI,
  output wire IRQ_P2F_CTI,
  output wire IRQ_P2F_GPIO,
  output wire IRQ_P2F_USB0,
  output wire IRQ_P2F_ENET0,
  output wire IRQ_P2F_ENET_WAKE0,
  output wire IRQ_P2F_SDIO0,
  output wire IRQ_P2F_I2C0,
  output wire IRQ_P2F_SPI0,
  output wire IRQ_P2F_UART0,
  output wire IRQ_P2F_CAN0,
  output wire IRQ_P2F_USB1,
  output wire IRQ_P2F_ENET1,
  output wire IRQ_P2F_ENET_WAKE1,
  output wire IRQ_P2F_SDIO1,
  output wire IRQ_P2F_I2C1,
  output wire IRQ_P2F_SPI1,
  output wire IRQ_P2F_UART1,
  output wire IRQ_P2F_CAN1,
  input  wire Core0_nFIQ,
  input  wire Core0_nIRQ,
  input  wire Core1_nFIQ,
  input  wire Core1_nIRQ,
  input  wire [15:0] IRQ_F2P,
  output wire EVENT_EVENTO,
  input wire EVENT_EVENTI,   
  output wire [1:0]  EVENT_STANDBYWFE,
  output wire [1:0]  EVENT_STANDBYWFI,  
   
  // Idle wire
  input wire FPGA_IDLE_n,
  
  // 4 fabric clks
  output wire FCLK0_CLK,
  output wire FCLK0_RESET_n,

  output wire FCLK1_CLK,
  output wire FCLK1_RESET_n,

  output wire FCLK2_CLK,
  output wire FCLK2_RESET_n,

  output wire FCLK3_CLK,
  output wire FCLK3_RESET_n,
  
  // PS Clock and Reset wires
  inout wire PS_SYSTEM_RESET,
  inout wire PS_CLK,         
  inout wire PS_POWER_ON_RESET,

  // DDR
  input [3:0] DDR_ARB,
  inout wire DDR_CAS_n,       
  inout wire DDR_CKE,         
  inout wire DDR_Clk_n,       
  inout wire DDR_Clk,         
  inout wire DDR_CS_n,         
  inout wire DDR_DRSTB,         
  inout wire DDR_ODT,         
  inout wire DDR_RAS_n,       
  inout wire DDR_WEB,
  inout wire [2:0]  DDR_BankAddr,      
  inout wire [14:0] DDR_Addr,          
  inout wire DDR_VRN,
  inout wire DDR_VRP,
  inout wire [3:0]  DDR_DM,            
  inout wire [31:0] DDR_DQ,          
  inout wire [3:0]  DDR_DQS_n,       
  inout wire [3:0]  DDR_DQS,         

  // AXI3+ (3 with some optional Axi4 wires)
  // direction is from PS point of view
  // 2 PS Master General Purpose ports
  // 2 PS Slave General Purpose ports
  // 1 PS Slave ACP port
  // 4 PS Slave High Performance ports

  //M_AXI_GP0
  output wire M_AXI_GP0_ARESET_n,
  output wire M_AXI_GP0_ARVALID,
  output wire M_AXI_GP0_AWVALID,
  output wire M_AXI_GP0_BREADY,
  output wire M_AXI_GP0_RREADY,
  output wire M_AXI_GP0_WLAST,
  output wire M_AXI_GP0_WVALID,
  output wire [11:0] M_AXI_GP0_ARID,
  output wire [11:0] M_AXI_GP0_AWID,
  output wire [11:0] M_AXI_GP0_WID,
  output wire [1:0] M_AXI_GP0_ARBURST,
  output wire [1:0] M_AXI_GP0_ARLOCK,
  output wire [1:0] M_AXI_GP0_ARSIZE,
  output wire [1:0] M_AXI_GP0_AWBURST,
  output wire [1:0] M_AXI_GP0_AWLOCK,
  output wire [1:0] M_AXI_GP0_AWSIZE,
  output wire [2:0] M_AXI_GP0_ARPROT,
  output wire [2:0] M_AXI_GP0_AWPROT,
  output wire [31:0] M_AXI_GP0_ARADDR,
  output wire [31:0] M_AXI_GP0_AWADDR,
  output wire [31:0] M_AXI_GP0_WDATA,
  output wire [3:0] M_AXI_GP0_ARCACHE,
  output wire [3:0] M_AXI_GP0_ARLEN,
  output wire [3:0] M_AXI_GP0_ARQOS,
  output wire [3:0] M_AXI_GP0_AWCACHE,
  output wire [3:0] M_AXI_GP0_AWLEN,
  output wire [3:0] M_AXI_GP0_AWQOS,
  output wire [3:0] M_AXI_GP0_WSTRB,
  input wire M_AXI_GP0_ACLK,
  input wire M_AXI_GP0_ARREADY,
  input wire M_AXI_GP0_AWREADY,
  input wire M_AXI_GP0_BVALID,
  input wire M_AXI_GP0_RLAST,
  input wire M_AXI_GP0_RVALID,
  input wire M_AXI_GP0_WREADY,
  input wire [11:0] M_AXI_GP0_BID,
  input wire [11:0] M_AXI_GP0_RID,
  input wire [1:0] M_AXI_GP0_BRESP,
  input wire [1:0] M_AXI_GP0_RRESP,
  input wire [31:0] M_AXI_GP0_RDATA,  

  //M_AXI_GP1
  output wire M_AXI_GP1_ARESET_n,
  output wire M_AXI_GP1_ARVALID,
  output wire M_AXI_GP1_AWVALID,
  output wire M_AXI_GP1_BREADY,
  output wire M_AXI_GP1_RREADY,
  output wire M_AXI_GP1_WLAST,
  output wire M_AXI_GP1_WVALID,
  output wire [11:0] M_AXI_GP1_ARID,
  output wire [11:0] M_AXI_GP1_AWID,
  output wire [11:0] M_AXI_GP1_WID,
  output wire [1:0] M_AXI_GP1_ARBURST,
  output wire [1:0] M_AXI_GP1_ARLOCK,
  output wire [1:0] M_AXI_GP1_ARSIZE,
  output wire [1:0] M_AXI_GP1_AWBURST,
  output wire [1:0] M_AXI_GP1_AWLOCK,
  output wire [1:0] M_AXI_GP1_AWSIZE,
  output wire [2:0] M_AXI_GP1_ARPROT,
  output wire [2:0] M_AXI_GP1_AWPROT,
  output wire [31:0] M_AXI_GP1_ARADDR,
  output wire [31:0] M_AXI_GP1_AWADDR,
  output wire [31:0] M_AXI_GP1_WDATA,
  output wire [3:0] M_AXI_GP1_ARCACHE,
  output wire [3:0] M_AXI_GP1_ARLEN,
  output wire [3:0] M_AXI_GP1_ARQOS,
  output wire [3:0] M_AXI_GP1_AWCACHE,
  output wire [3:0] M_AXI_GP1_AWLEN,
  output wire [3:0] M_AXI_GP1_AWQOS,
  output wire [3:0] M_AXI_GP1_WSTRB,
  input wire M_AXI_GP1_ACLK,
  input wire M_AXI_GP1_ARREADY,
  input wire M_AXI_GP1_AWREADY,
  input wire M_AXI_GP1_BVALID,
  input wire M_AXI_GP1_RLAST,
  input wire M_AXI_GP1_RVALID,
  input wire M_AXI_GP1_WREADY,  
  input wire [11:0] M_AXI_GP1_BID,
  input wire [11:0] M_AXI_GP1_RID,
  input wire [1:0] M_AXI_GP1_BRESP,
  input wire [1:0] M_AXI_GP1_RRESP,
  input wire [31:0] M_AXI_GP1_RDATA,
  
  // S_AXI_GP0
  output wire S_AXI_GP0_ARESET_n,
  output wire S_AXI_GP0_ARREADY,
  output wire S_AXI_GP0_AWREADY,
  output wire S_AXI_GP0_BVALID,
  output wire S_AXI_GP0_RLAST,
  output wire S_AXI_GP0_RVALID,
  output wire S_AXI_GP0_WREADY,  
  output wire [1:0] S_AXI_GP0_BRESP,
  output wire [1:0] S_AXI_GP0_RRESP,
  output wire [31:0] S_AXI_GP0_RDATA,
  output wire [5:0] S_AXI_GP0_BID,
  output wire [5:0] S_AXI_GP0_RID,
  input wire S_AXI_GP0_ACLK,
  input wire S_AXI_GP0_ARVALID,
  input wire S_AXI_GP0_AWVALID,
  input wire S_AXI_GP0_BREADY,
  input wire S_AXI_GP0_RREADY,
  input wire S_AXI_GP0_WLAST,
  input wire S_AXI_GP0_WVALID,
  input wire [1:0] S_AXI_GP0_ARBURST,
  input wire [1:0] S_AXI_GP0_ARLOCK,
  input wire [1:0] S_AXI_GP0_ARSIZE,
  input wire [1:0] S_AXI_GP0_AWBURST,
  input wire [1:0] S_AXI_GP0_AWLOCK,
  input wire [1:0] S_AXI_GP0_AWSIZE,
  input wire [2:0] S_AXI_GP0_ARPROT,
  input wire [2:0] S_AXI_GP0_AWPROT,
  input wire [31:0] S_AXI_GP0_ARADDR,
  input wire [31:0] S_AXI_GP0_AWADDR,
  input wire [31:0] S_AXI_GP0_WDATA,
  input wire [3:0] S_AXI_GP0_ARCACHE,
  input wire [3:0] S_AXI_GP0_ARLEN,
  input wire [3:0] S_AXI_GP0_ARQOS,
  input wire [3:0] S_AXI_GP0_AWCACHE,
  input wire [3:0] S_AXI_GP0_AWLEN,
  input wire [3:0] S_AXI_GP0_AWQOS,
  input wire [3:0] S_AXI_GP0_WSTRB,
  input wire [5:0] S_AXI_GP0_ARID,
  input wire [5:0] S_AXI_GP0_AWID,
  input wire [5:0] S_AXI_GP0_WID,  

  // S_AXI_GP1
  output wire S_AXI_GP1_ARESET_n,
  output wire S_AXI_GP1_ARREADY,
  output wire S_AXI_GP1_AWREADY,
  output wire S_AXI_GP1_BVALID,
  output wire S_AXI_GP1_RLAST,
  output wire S_AXI_GP1_RVALID,
  output wire S_AXI_GP1_WREADY,  
  output wire [1:0] S_AXI_GP1_BRESP,
  output wire [1:0] S_AXI_GP1_RRESP,
  output wire [31:0] S_AXI_GP1_RDATA,
  output wire [5:0] S_AXI_GP1_BID,
  output wire [5:0] S_AXI_GP1_RID,
  input wire S_AXI_GP1_ACLK,
  input wire S_AXI_GP1_ARVALID,
  input wire S_AXI_GP1_AWVALID,
  input wire S_AXI_GP1_BREADY,
  input wire S_AXI_GP1_RREADY,
  input wire S_AXI_GP1_WLAST,
  input wire S_AXI_GP1_WVALID,
  input wire [1:0] S_AXI_GP1_ARBURST,
  input wire [1:0] S_AXI_GP1_ARLOCK,
  input wire [1:0] S_AXI_GP1_ARSIZE,
  input wire [1:0] S_AXI_GP1_AWBURST,
  input wire [1:0] S_AXI_GP1_AWLOCK,
  input wire [1:0] S_AXI_GP1_AWSIZE,
  input wire [2:0] S_AXI_GP1_ARPROT,
  input wire [2:0] S_AXI_GP1_AWPROT,
  input wire [31:0] S_AXI_GP1_ARADDR,
  input wire [31:0] S_AXI_GP1_AWADDR,
  input wire [31:0] S_AXI_GP1_WDATA,
  input wire [3:0] S_AXI_GP1_ARCACHE,
  input wire [3:0] S_AXI_GP1_ARLEN,
  input wire [3:0] S_AXI_GP1_ARQOS,
  input wire [3:0] S_AXI_GP1_AWCACHE,
  input wire [3:0] S_AXI_GP1_AWLEN,
  input wire [3:0] S_AXI_GP1_AWQOS,
  input wire [3:0] S_AXI_GP1_WSTRB,
  input wire [5:0] S_AXI_GP1_ARID,
  input wire [5:0] S_AXI_GP1_AWID,
  input wire [5:0] S_AXI_GP1_WID, 

  //S_AXI_ACP
  output wire S_AXI_ACP_ARESET_n,
  output wire S_AXI_ACP_ARREADY,
  output wire S_AXI_ACP_AWREADY,
  output wire S_AXI_ACP_BVALID,
  output wire S_AXI_ACP_RLAST,
  output wire S_AXI_ACP_RVALID,
  output wire S_AXI_ACP_WREADY,  
  output wire [1:0] S_AXI_ACP_BRESP,
  output wire [1:0] S_AXI_ACP_RRESP,
  output wire [2 : 0] S_AXI_ACP_BID,
  output wire [2 : 0] S_AXI_ACP_RID,
  output wire [63:0] S_AXI_ACP_RDATA,
  input wire S_AXI_ACP_ACLK,
  input wire S_AXI_ACP_ARVALID,
  input wire S_AXI_ACP_AWVALID,
  input wire S_AXI_ACP_BREADY,
  input wire S_AXI_ACP_RREADY,
  input wire S_AXI_ACP_WLAST,
  input wire S_AXI_ACP_WVALID,
  input wire [2:0] S_AXI_ACP_ARID,
  input wire [2:0] S_AXI_ACP_ARPROT,
  input wire [2:0] S_AXI_ACP_AWID,
  input wire [2:0] S_AXI_ACP_AWPROT,
  input wire [2:0] S_AXI_ACP_WID,
  input wire [31:0] S_AXI_ACP_ARADDR,
  input wire [31:0] S_AXI_ACP_AWADDR,
  input wire [3:0] S_AXI_ACP_ARCACHE,
  input wire [3:0] S_AXI_ACP_ARLEN,
  input wire [3:0] S_AXI_ACP_ARQOS,
  input wire [3:0] S_AXI_ACP_AWCACHE,
  input wire [3:0] S_AXI_ACP_AWLEN,
  input wire [3:0] S_AXI_ACP_AWQOS,
  input wire [1:0] S_AXI_ACP_ARBURST,
  input wire [1:0] S_AXI_ACP_ARLOCK,
  input wire [1:0] S_AXI_ACP_ARSIZE,
  input wire [1:0] S_AXI_ACP_AWBURST,
  input wire [1:0] S_AXI_ACP_AWLOCK,
  input wire [1:0] S_AXI_ACP_AWSIZE,
  input wire [4:0] S_AXI_ACP_ARUSER,
  input wire [4:0] S_AXI_ACP_AWUSER,
  input wire [63:0] S_AXI_ACP_WDATA,
  input wire [7:0] S_AXI_ACP_WSTRB, 

  // AXI HP0
  output wire S_AXI_HP0_ARESET_n,
  output wire S_AXI_HP0_ARREADY,
  output wire S_AXI_HP0_AWREADY,
  output wire S_AXI_HP0_BVALID,
  output wire S_AXI_HP0_RLAST,
  output wire S_AXI_HP0_RVALID,
  output wire S_AXI_HP0_WREADY,  
  output wire [1:0] S_AXI_HP0_BRESP,
  output wire [1:0] S_AXI_HP0_RRESP,
  output wire [5:0] S_AXI_HP0_BID,
  output wire [5:0] S_AXI_HP0_RID,
  output wire [63:0] S_AXI_HP0_RDATA,
  output wire [7:0] S_AXI_HP0_RCOUNT,
  output wire [7:0] S_AXI_HP0_WCOUNT,
  output wire [2:0] S_AXI_HP0_RACOUNT,
  output wire [5:0] S_AXI_HP0_WACOUNT,
  input wire S_AXI_HP0_ACLK,
  input wire S_AXI_HP0_ARVALID,
  input wire S_AXI_HP0_AWVALID,
  input wire S_AXI_HP0_BREADY,
  input wire S_AXI_HP0_RDISSUECAP1_EN,
  input wire S_AXI_HP0_RREADY,
  input wire S_AXI_HP0_WLAST,
  input wire S_AXI_HP0_WRISSUECAP1_EN,
  input wire S_AXI_HP0_WVALID,
  input wire [1:0] S_AXI_HP0_ARBURST,
  input wire [1:0] S_AXI_HP0_ARLOCK,
  input wire [1:0] S_AXI_HP0_ARSIZE,
  input wire [1:0] S_AXI_HP0_AWBURST,
  input wire [1:0] S_AXI_HP0_AWLOCK,
  input wire [1:0] S_AXI_HP0_AWSIZE,
  input wire [2:0] S_AXI_HP0_ARPROT,
  input wire [2:0] S_AXI_HP0_AWPROT,
  input wire [31:0] S_AXI_HP0_ARADDR,
  input wire [31:0] S_AXI_HP0_AWADDR,
  input wire [3:0] S_AXI_HP0_ARCACHE,
  input wire [3:0] S_AXI_HP0_ARLEN,
  input wire [3:0] S_AXI_HP0_ARQOS,
  input wire [3:0] S_AXI_HP0_AWCACHE,
  input wire [3:0] S_AXI_HP0_AWLEN,
  input wire [3:0] S_AXI_HP0_AWQOS,
  input wire [5:0] S_AXI_HP0_ARID,
  input wire [5:0] S_AXI_HP0_AWID,
  input wire [5:0] S_AXI_HP0_WID,
  input wire [63:0] S_AXI_HP0_WDATA,
  input wire [7:0] S_AXI_HP0_WSTRB,

  // AXI HP1
  output wire S_AXI_HP1_ARESET_n,
  output wire S_AXI_HP1_ARREADY,
  output wire S_AXI_HP1_AWREADY,
  output wire S_AXI_HP1_BVALID,
  output wire S_AXI_HP1_RLAST,
  output wire S_AXI_HP1_RVALID,
  output wire S_AXI_HP1_WREADY,  
  output wire [1:0] S_AXI_HP1_BRESP,
  output wire [1:0] S_AXI_HP1_RRESP,
  output wire [5:0] S_AXI_HP1_BID,
  output wire [5:0] S_AXI_HP1_RID,
  output wire [63:0] S_AXI_HP1_RDATA,
  output wire [7:0] S_AXI_HP1_RCOUNT,
  output wire [7:0] S_AXI_HP1_WCOUNT,
  output wire [2:0] S_AXI_HP1_RACOUNT,
  output wire [5:0] S_AXI_HP1_WACOUNT,
  input wire S_AXI_HP1_ACLK,
  input wire S_AXI_HP1_ARVALID,
  input wire S_AXI_HP1_AWVALID,
  input wire S_AXI_HP1_BREADY,
  input wire S_AXI_HP1_RDISSUECAP1_EN,
  input wire S_AXI_HP1_RREADY,
  input wire S_AXI_HP1_WLAST,
  input wire S_AXI_HP1_WRISSUECAP1_EN,
  input wire S_AXI_HP1_WVALID,
  input wire [1:0] S_AXI_HP1_ARBURST,
  input wire [1:0] S_AXI_HP1_ARLOCK,
  input wire [1:0] S_AXI_HP1_ARSIZE,
  input wire [1:0] S_AXI_HP1_AWBURST,
  input wire [1:0] S_AXI_HP1_AWLOCK,
  input wire [1:0] S_AXI_HP1_AWSIZE,
  input wire [2:0] S_AXI_HP1_ARPROT,
  input wire [2:0] S_AXI_HP1_AWPROT,
  input wire [31:0] S_AXI_HP1_ARADDR,
  input wire [31:0] S_AXI_HP1_AWADDR,
  input wire [3:0] S_AXI_HP1_ARCACHE,
  input wire [3:0] S_AXI_HP1_ARLEN,
  input wire [3:0] S_AXI_HP1_ARQOS,
  input wire [3:0] S_AXI_HP1_AWCACHE,
  input wire [3:0] S_AXI_HP1_AWLEN,
  input wire [3:0] S_AXI_HP1_AWQOS,
  input wire [5:0] S_AXI_HP1_ARID,
  input wire [5:0] S_AXI_HP1_AWID,
  input wire [5:0] S_AXI_HP1_WID,
  input wire [63:0] S_AXI_HP1_WDATA,
  input wire [7:0] S_AXI_HP1_WSTRB,

  // S_AXI_HP2
  output wire S_AXI_HP2_ARESET_n,
  output wire S_AXI_HP2_ARREADY,
  output wire S_AXI_HP2_AWREADY,
  output wire S_AXI_HP2_BVALID,
  output wire S_AXI_HP2_RLAST,
  output wire S_AXI_HP2_RVALID,
  output wire S_AXI_HP2_WREADY,  
  output wire [1:0] S_AXI_HP2_BRESP,
  output wire [1:0] S_AXI_HP2_RRESP,
  output wire [5:0] S_AXI_HP2_BID,
  output wire [5:0] S_AXI_HP2_RID,
  output wire [63:0] S_AXI_HP2_RDATA,
  output wire [7:0] S_AXI_HP2_RCOUNT,
  output wire [7:0] S_AXI_HP2_WCOUNT,
  output wire [2:0] S_AXI_HP2_RACOUNT,
  output wire [5:0] S_AXI_HP2_WACOUNT,
  input wire S_AXI_HP2_ACLK,
  input wire S_AXI_HP2_ARVALID,
  input wire S_AXI_HP2_AWVALID,
  input wire S_AXI_HP2_BREADY,
  input wire S_AXI_HP2_RDISSUECAP1_EN,
  input wire S_AXI_HP2_RREADY,
  input wire S_AXI_HP2_WLAST,
  input wire S_AXI_HP2_WRISSUECAP1_EN,
  input wire S_AXI_HP2_WVALID,
  input wire [1:0] S_AXI_HP2_ARBURST,
  input wire [1:0] S_AXI_HP2_ARLOCK,
  input wire [1:0] S_AXI_HP2_ARSIZE,
  input wire [1:0] S_AXI_HP2_AWBURST,
  input wire [1:0] S_AXI_HP2_AWLOCK,
  input wire [1:0] S_AXI_HP2_AWSIZE,
  input wire [2:0] S_AXI_HP2_ARPROT,
  input wire [2:0] S_AXI_HP2_AWPROT,
  input wire [31:0] S_AXI_HP2_ARADDR,
  input wire [31:0] S_AXI_HP2_AWADDR,
  input wire [3:0] S_AXI_HP2_ARCACHE,
  input wire [3:0] S_AXI_HP2_ARLEN,
  input wire [3:0] S_AXI_HP2_ARQOS,
  input wire [3:0] S_AXI_HP2_AWCACHE,
  input wire [3:0] S_AXI_HP2_AWLEN,
  input wire [3:0] S_AXI_HP2_AWQOS,
  input wire [5:0] S_AXI_HP2_ARID,
  input wire [5:0] S_AXI_HP2_AWID,
  input wire [5:0] S_AXI_HP2_WID,
  input wire [63:0] S_AXI_HP2_WDATA,
  input wire [7:0] S_AXI_HP2_WSTRB,

  // S_AXI_HP_3
  output wire S_AXI_HP3_ARESET_n,
  output wire S_AXI_HP3_ARREADY,
  output wire S_AXI_HP3_AWREADY,
  output wire S_AXI_HP3_BVALID,
  output wire S_AXI_HP3_RLAST,
  output wire S_AXI_HP3_RVALID,
  output wire S_AXI_HP3_WREADY,  
  output wire [1:0] S_AXI_HP3_BRESP,
  output wire [1:0] S_AXI_HP3_RRESP,
  output wire [5:0] S_AXI_HP3_BID,
  output wire [5:0] S_AXI_HP3_RID,
  output wire [63:0] S_AXI_HP3_RDATA,
  output wire [7:0] S_AXI_HP3_RCOUNT,
  output wire [7:0] S_AXI_HP3_WCOUNT,
  output wire [2:0] S_AXI_HP3_RACOUNT,
  output wire [5:0] S_AXI_HP3_WACOUNT,
  input wire S_AXI_HP3_ACLK,
  input wire S_AXI_HP3_ARVALID,
  input wire S_AXI_HP3_AWVALID,
  input wire S_AXI_HP3_BREADY,
  input wire S_AXI_HP3_RDISSUECAP1_EN,
  input wire S_AXI_HP3_RREADY,
  input wire S_AXI_HP3_WLAST,
  input wire S_AXI_HP3_WRISSUECAP1_EN,
  input wire S_AXI_HP3_WVALID,
  input wire [1:0] S_AXI_HP3_ARBURST,
  input wire [1:0] S_AXI_HP3_ARLOCK,
  input wire [1:0] S_AXI_HP3_ARSIZE,
  input wire [1:0] S_AXI_HP3_AWBURST,
  input wire [1:0] S_AXI_HP3_AWLOCK,
  input wire [1:0] S_AXI_HP3_AWSIZE,
  input wire [2:0] S_AXI_HP3_ARPROT,
  input wire [2:0] S_AXI_HP3_AWPROT,
  input wire [31:0] S_AXI_HP3_ARADDR,
  input wire [31:0] S_AXI_HP3_AWADDR,
  input wire [3:0] S_AXI_HP3_ARCACHE,
  input wire [3:0] S_AXI_HP3_ARLEN,
  input wire [3:0] S_AXI_HP3_ARQOS,
  input wire [3:0] S_AXI_HP3_AWCACHE,
  input wire [3:0] S_AXI_HP3_AWLEN,
  input wire [3:0] S_AXI_HP3_AWQOS,
  input wire [5:0] S_AXI_HP3_ARID,
  input wire [5:0] S_AXI_HP3_AWID,
  input wire [5:0] S_AXI_HP3_WID,
  input wire [63:0] S_AXI_HP3_WDATA,
  input wire [7:0] S_AXI_HP3_WSTRB

);

  PS7 PS7_i (
    // 2x CAN
	  .EMIOCAN0PHYTX	          (CAN0_PHY_TX),
	  .EMIOCAN0PHYRX	          (CAN0_PHY_RX),
	  .EMIOCAN1PHYTX	          (CAN1_PHY_TX),
	  .EMIOCAN1PHYRX	          (CAN1_PHY_RX),

    // 2x gigabit ethernet
	  .EMIOENET0EXTINTIN        (ENET0_EXT_INTIN),  
	  .EMIOENET0GMIICOL         (ENET0_GMII_COL),
	  .EMIOENET0GMIICRS         (ENET0_GMII_CRS),
	  .EMIOENET0GMIIRXCLK       (ENET0_GMII_RX_CLK),
	  .EMIOENET0GMIIRXD         (ENET0_GMII_RXD),
	  .EMIOENET0GMIIRXDV        (ENET0_GMII_RX_DV),
	  .EMIOENET0GMIIRXER        (ENET0_GMII_RX_ER),
	  .EMIOENET0GMIITXCLK       (ENET0_GMII_TX_CLK),
	  .EMIOENET0MDIOI           (ENET0_MDIO_I),
	  .EMIOENET0GMIITXD	        (ENET0_GMII_TXD),
    .EMIOENET0GMIITXEN	      (ENET0_GMII_TX_EN),
	  .EMIOENET0GMIITXER        (ENET0_GMII_TX_ER), 
	  .EMIOENET0MDIOMDC	        (ENET0_MDIO_MDC),
	  .EMIOENET0MDIOO	          (ENET0_MDIO_O),
	  .EMIOENET0MDIOTN	        (ENET0_MDIO_T_n),
	  .EMIOENET0PTPDELAYREQRX   (ENET0_PTP_DELAY_REQ_RX),
	  .EMIOENET0PTPDELAYREQTX   (ENET0_PTP_DELAY_REQ_TX),
	  .EMIOENET0PTPPDELAYREQRX  (ENET0_PTP_PDELAY_REQ_RX),
	  .EMIOENET0PTPPDELAYREQTX  (ENET0_PTP_PDELAY_REQ_TX),
	  .EMIOENET0PTPPDELAYRESPRX (ENET0_PTP_PDELAY_RESP_RX),
	  .EMIOENET0PTPPDELAYRESPTX (ENET0_PTP_PDELAY_RESP_TX),
	  .EMIOENET0PTPSYNCFRAMERX  (ENET0_PTP_SYNC_FRAME_RX),
	  .EMIOENET0PTPSYNCFRAMETX  (ENET0_PTP_SYNC_FRAME_TX),
	  .EMIOENET0SOFRX           (ENET0_SOF_RX),
	  .EMIOENET0SOFTX           (ENET0_SOF_TX),

	  .EMIOENET1EXTINTIN        (ENET1_EXT_INTIN),    
	  .EMIOENET1GMIICOL         (ENET1_GMII_COL),
	  .EMIOENET1GMIICRS         (ENET1_GMII_CRS),
	  .EMIOENET1GMIIRXCLK       (ENET1_GMII_RX_CLK),
	  .EMIOENET1GMIIRXD         (ENET1_GMII_RXD),
	  .EMIOENET1GMIIRXDV        (ENET1_GMII_RX_DV),
	  .EMIOENET1GMIIRXER        (ENET1_GMII_RX_ER),
	  .EMIOENET1GMIITXCLK       (ENET1_GMII_TX_CLK),
	  .EMIOENET1MDIOI           (ENET1_MDIO_I),
	  .EMIOENET1GMIITXD	        (ENET1_GMII_TXD),
	  .EMIOENET1GMIITXEN	      (ENET1_GMII_TX_EN),
	  .EMIOENET1GMIITXER	      (ENET1_GMII_TX_ER),
	  .EMIOENET1MDIOMDC	        (ENET1_MDIO_MDC),
	  .EMIOENET1MDIOO	          (ENET1_MDIO_O),
	  .EMIOENET1MDIOTN	        (ENET1_MDIO_T_n),
	  .EMIOENET1PTPDELAYREQRX   (ENET1_PTP_DELAY_REQ_RX),
	  .EMIOENET1PTPDELAYREQTX   (ENET1_PTP_DELAY_REQ_TX),
	  .EMIOENET1PTPPDELAYREQRX  (ENET1_PTP_PDELAY_REQ_RX),
	  .EMIOENET1PTPPDELAYREQTX  (ENET1_PTP_PDELAY_REQ_TX),
	  .EMIOENET1PTPPDELAYRESPRX (ENET1_PTP_PDELAY_RESP_RX),
	  .EMIOENET1PTPPDELAYRESPTX (ENET1_PTP_PDELAY_RESP_TX),
	  .EMIOENET1PTPSYNCFRAMERX  (ENET1_PTP_SYNC_FRAME_RX),
	  .EMIOENET1PTPSYNCFRAMETX  (ENET1_PTP_SYNC_FRAME_TX),
	  .EMIOENET1SOFRX           (ENET1_SOF_RX),
	  .EMIOENET1SOFTX           (ENET1_SOF_TX),

    // 4x DMA
	  .DMA0ACLK		              (DMA0_ACLK),
	  .DMA0RSTN		              (DMA0_RESET_n),  
	  .DMA0DATYPE		            (DMA0_DATYPE),
	  .DMA0DAVALID		          (DMA0_DAVALID),
	  .DMA0DRREADY		          (DMA0_DRREADY),  
	  .DMA0DAREADY		          (DMA0_DAREADY),
	  .DMA0DRLAST		            (DMA0_DRLAST),
	  .DMA0DRTYPE               (DMA0_DRTYPE),
	  .DMA0DRVALID		          (DMA0_DRVALID),

	  .DMA1ACLK		              (DMA1_ACLK),
	  .DMA1RSTN		              (DMA1_RESET_n),
	  .DMA1DATYPE		            (DMA1_DATYPE),
	  .DMA1DAVALID		          (DMA1_DAVALID),
	  .DMA1DRREADY		          (DMA1_DRREADY),
	  .DMA1DAREADY		          (DMA1_DAREADY),
	  .DMA1DRLAST		            (DMA1_DRLAST),
	  .DMA1DRTYPE               (DMA1_DRTYPE),  
	  .DMA1DRVALID		          (DMA1_DRVALID),

	  .DMA2ACLK		              (DMA2_ACLK),
	  .DMA2RSTN		              (DMA2_RESET_n),
	  .DMA2DATYPE		            (DMA2_DATYPE),
	  .DMA2DAVALID		          (DMA2_DAVALID),
	  .DMA2DRREADY		          (DMA2_DRREADY),
	  .DMA2DAREADY		          (DMA2_DAREADY),
	  .DMA2DRLAST		            (DMA2_DRLAST),
	  .DMA2DRTYPE               (DMA2_DRTYPE),    
	  .DMA2DRVALID		          (DMA2_DRVALID),

	  .DMA3ACLK		              (DMA3_ACLK),
	  .DMA3RSTN		              (DMA3_RESET_n),
	  .DMA3DAREADY		          (DMA3_DAREADY),
	  .DMA3DRLAST		            (DMA3_DRLAST),
	  .DMA3DRTYPE               (DMA3_DRTYPE),
	  .DMA3DRVALID		          (DMA3_DRVALID),
	  .DMA3DATYPE		            (DMA3_DATYPE),
	  .DMA3DAVALID		          (DMA3_DAVALID),
	  .DMA3DRREADY		          (DMA3_DRREADY),

    // gpio 
	  .EMIOGPIOI	              (GPIO_I),
	  .EMIOGPIOO	              (GPIO_O),
	  .EMIOGPIOTN	              (GPIO_T_n),
	  .MIO			                (MIO),
	  
    // 2x I2C
    .EMIOI2C0SCLO             (I2C0_SCL_O),
	  .EMIOI2C0SCLTN            (I2C0_SCL_T_n),
	  .EMIOI2C0SDAO	            (I2C0_SDA_O),
	  .EMIOI2C0SDATN	          (I2C0_SDA_T_n),
	  .EMIOI2C0SCLI	            (I2C0_SCL_I),
	  .EMIOI2C0SDAI	            (I2C0_SDA_I),

	  .EMIOI2C1SCLO	            (I2C1_SCL_O),
	  .EMIOI2C1SCLTN            (I2C1_SCL_T_n),
	  .EMIOI2C1SDAO	            (I2C1_SDA_O),
	  .EMIOI2C1SDATN	          (I2C1_SDA_T_n),
	  .EMIOI2C1SCLI	            (I2C1_SCL_I),
	  .EMIOI2C1SDAI	            (I2C1_SDA_I),

	  
    // 2x SDIO
	  .EMIOSDIO0BUSPOW          (SDIO0_BUSPOW),  
    .EMIOSDIO0CLK		          (SDIO0_CLK),
	  .EMIOSDIO0CMDO	          (SDIO0_CMD_O),
	  .EMIOSDIO0CMDTN	          (SDIO0_CMD_T_n),
	  .EMIOSDIO0DATAO	          (SDIO0_DATA_O),
	  .EMIOSDIO0DATATN	        (SDIO0_DATA_T_n),
	  .EMIOSDIO0LED             (SDIO0_LED),
	  .EMIOSDIO0BUSVOLT         (SDIO0_BUSVOLT), 
	  .EMIOSDIO0CDN             (SDIO0_CDN),
	  .EMIOSDIO0CLKFB	          (SDIO0_CLK_FB),
	  .EMIOSDIO0CMDI	          (SDIO0_CMD_I),
	  .EMIOSDIO0DATAI	          (SDIO0_DATA_I),
	  .EMIOSDIO0WP              (SDIO0_WP),

	  .EMIOSDIO1BUSPOW          (SDIO1_BUSPOW),  
	  .EMIOSDIO1CLK             (SDIO1_CLK),
	  .EMIOSDIO1CMDO            (SDIO1_CMD_O),
	  .EMIOSDIO1CMDTN           (SDIO1_CMD_T_n),
	  .EMIOSDIO1DATAO           (SDIO1_DATA_O),
	  .EMIOSDIO1DATATN          (SDIO1_DATA_T_n),
	  .EMIOSDIO1LED             (SDIO1_LED),
	  .EMIOSDIO1CDN             (SDIO1_CDN),
	  .EMIOSDIO1CLKFB	          (SDIO1_CLK_FB),
	  .EMIOSDIO1CMDI	          (SDIO1_CMD_I),
	  .EMIOSDIO1DATAI	          (SDIO1_DATA_I),
	  .EMIOSDIO1WP              (SDIO1_WP),
	  .EMIOSDIO1BUSVOLT         (SDIO1_BUSVOLT),  

    // 2x SPI
	  .EMIOSPI0MO		            (SPI0_MOSI_O),
	  .EMIOSPI0MOTN	            (SPI0_MOSI_T_n),
	  .EMIOSPI0SCLKO	          (SPI0_SCLK_O),
	  .EMIOSPI0SCLKTN	          (SPI0_SCLK_T_n),
	  .EMIOSPI0SO		            (SPI0_MISO_O),
	  .EMIOSPI0STN	            (SPI0_MISO_T_n),
	  .EMIOSPI0SSON	            ({SPI0_SS2_O,SPI0_SS1_O,SPI0_SS_O}),
	  .EMIOSPI0SSNTN	          (SPI0_SS_T_n),
	  .EMIOSPI0MI		            (SPI0_MISO_I),
	  .EMIOSPI0SCLKI	          (SPI0_SCLK_I),
	  .EMIOSPI0SI		            (SPI0_MOSI_I),
	  .EMIOSPI0SSIN 	          (SPI0_SS_I),

	  .EMIOSPI1MO		            (SPI1_MOSI_O),
	  .EMIOSPI1MOTN	            (SPI1_MOSI_T_n),
	  .EMIOSPI1SCLKO	          (SPI1_SCLK_O),
	  .EMIOSPI1SCLKTN	          (SPI1_SCLK_T_n),
	  .EMIOSPI1SO		            (SPI1_MISO_O),
	  .EMIOSPI1STN	            (SPI1_MISO_T_n),
	  .EMIOSPI1SSON	            ({SPI1_SS2_O,SPI1_SS1_O,SPI1_SS_O}),
	  .EMIOSPI1SSNTN	          (SPI1_SS_T_n),
	  .EMIOSPI1MI		            (SPI1_MISO_I),
	  .EMIOSPI1SCLKI	          (SPI1_SCLK_I),
	  .EMIOSPI1SI		            (SPI1_MOSI_I),
	  .EMIOSPI1SSIN	            (SPI1_SS_I),

    // jtag, trace and debug
	  .EMIOTRACECLK		          (TRACE_CLK),
	  .EMIOTRACECTL		          (TRACE_CTL),
	  .EMIOTRACEDATA	          (TRACE_DATA),
	  .EMIOTTC0CLKI	            ({TTC0_CLK2_IN, TTC0_CLK1_IN, TTC0_CLK0_IN}),
	  .EMIOTTC0WAVEO	          ({TTC0_WAVE2_OUT,TTC0_WAVE1_OUT,TTC0_WAVE0_OUT}),
	  .EMIOTTC1CLKI	            ({TTC1_CLK2_IN, TTC1_CLK1_IN, TTC1_CLK0_IN}),
	  .EMIOTTC1WAVEO	          ({TTC1_WAVE2_OUT,TTC1_WAVE1_OUT,TTC1_WAVE0_OUT}),

	  .FTMDTRACEINCLOCK	        (FTMD_TRACEIN_CLK ),
	  .FTMDTRACEINATID	        (FTMD_TRACEIN_ATID),  
	  .FTMDTRACEINDATA	        (FTMD_TRACEIN_DATA),
	  .FTMDTRACEINVALID	        (FTMD_TRACEIN_VALID),

	  .FTMTP2FDEBUG		          (FTMT_P2F_DEBUG),
	  .FTMTP2FTRIG		          ({FTMT_P2F_TRIG_3,FTMT_P2F_TRIG_2,FTMT_P2F_TRIG_1,FTMT_P2F_TRIG_0}),
	  .FTMTP2FTRIGACK	          ({FTMT_P2F_TRIGACK_3,FTMT_P2F_TRIGACK_2,FTMT_P2F_TRIGACK_1,FTMT_P2F_TRIGACK_0}),  

	  .FTMTF2PDEBUG		          (FTMT_F2P_DEBUG),
	  .FTMTF2PTRIG		          ({FTMT_F2P_TRIG_3,FTMT_F2P_TRIG_2,FTMT_F2P_TRIG_1,FTMT_F2P_TRIG_0}),
	  .FTMTF2PTRIGACK	          ({FTMT_F2P_TRIGACK_3,FTMT_F2P_TRIGACK_2,FTMT_F2P_TRIGACK_1,FTMT_F2P_TRIGACK_0}),

    .EMIOPJTAGTDO  	          (PJTAG_TDO_O),
	  .EMIOPJTAGTDTN	          (PJTAG_TDO_T_n),
	  .EMIOPJTAGTCK		          (PJTAG_TCK),
	  .EMIOPJTAGTDI		          (PJTAG_TDI),
	  .EMIOPJTAGTMS		          (PJTAG_TMS),

    // 2xUART
    .EMIOUART0DTRN	          (UART0_DTRN),
	  .EMIOUART0RTSN	          (UART0_RTSN),
	  .EMIOUART0TX		          (UART0_TX),
	  .EMIOUART0CTSN	          (UART0_CTSN),
	  .EMIOUART0DCDN	          (UART0_DCDN),
	  .EMIOUART0DSRN	          (UART0_DSRN),
	  .EMIOUART0RIN		          (UART0_RIN),
	  .EMIOUART0RX		          (UART0_RX),

	  .EMIOUART1DTRN	          (UART1_DTRN),
	  .EMIOUART1RTSN	          (UART1_RTSN),
	  .EMIOUART1TX		          (UART1_TX),
	  .EMIOUART1CTSN	          (UART1_CTSN),
	  .EMIOUART1DCDN	          (UART1_DCDN),
	  .EMIOUART1DSRN	          (UART1_DSRN),
	  .EMIOUART1RIN		          (UART1_RIN),
	  .EMIOUART1RX		          (UART1_RX),

    // Misc
	  .PSCLK		                (PS_CLK),
	  .PSPORB		                (PS_POWER_ON_RESET),
	  .PSSRSTB		              (PS_SYSTEM_RESET),
	  .FPGAIDLEN		            (FPGA_IDLE_n),
	  .EMIOSRAMINTIN            (SRAM_INTIN),

    // 2x USB 
	  .EMIOUSB0PORTINDCTL       (USB0_PORT_INDCTL),  
	  .EMIOUSB0VBUSPWRSELECT    (USB0_VBUS_PWRSELECT),
	  .EMIOUSB0VBUSPWRFAULT     (USB0_VBUS_PWRFAULT),
	  .EMIOUSB1PORTINDCTL       (USB1_PORT_INDCTL),
	  .EMIOUSB1VBUSPWRSELECT    (USB1_VBUS_PWRSELECT),  
	  .EMIOUSB1VBUSPWRFAULT     (USB1_VBUS_PWRFAULT),  

    // Watch Dog
	  .EMIOWDTRSTO    	        (WDT_RST_OUT),
	  .EMIOWDTCLKI		          (WDT_CLK_IN),  

    // events and interrupts
	  .EVENTEVENTO              (EVENT_EVENTO),
	  .EVENTSTANDBYWFE          (EVENT_STANDBYWFE),
	  .EVENTSTANDBYWFI          (EVENT_STANDBYWFI),  
	  .IRQP2F		                ({IRQ_P2F_DMAC_ABORT, IRQ_P2F_DMAC7, IRQ_P2F_DMAC6, IRQ_P2F_DMAC5, IRQ_P2F_DMAC4, IRQ_P2F_DMAC3, IRQ_P2F_DMAC2, IRQ_P2F_DMAC1, IRQ_P2F_DMAC0, IRQ_P2F_SMC, IRQ_P2F_QSPI, IRQ_P2F_CTI, IRQ_P2F_GPIO, IRQ_P2F_USB0, IRQ_P2F_ENET0, IRQ_P2F_ENET_WAKE0, IRQ_P2F_SDIO0, IRQ_P2F_I2C0, IRQ_P2F_SPI0, IRQ_P2F_UART0, IRQ_P2F_CAN0, IRQ_P2F_USB1, IRQ_P2F_ENET1, IRQ_P2F_ENET_WAKE1, IRQ_P2F_SDIO1, IRQ_P2F_I2C1, IRQ_P2F_SPI1, IRQ_P2F_UART1, IRQ_P2F_CAN1}),    
	  .EVENTEVENTI              (EVENT_EVENTI),
	  .IRQF2P		                ({Core1_nFIQ,Core0_nFIQ,Core1_nIRQ,Core0_nIRQ,IRQ_F2P[15:0]}),  

    // 4 x FCLK
	  .FCLKCLK		              ({FCLK3_CLK, FCLK2_CLK, FCLK1_CLK, FCLK0_CLK}),
 	  .FCLKRESETN		            ({FCLK3_RESET_n,FCLK2_RESET_n,FCLK1_RESET_n,FCLK0_RESET_n}),
	  .FCLKCLKTRIGN		          ({'b0, 'b0, 'b0, 'b0}),

    // DDR
    .DDRARB                   (DDR_ARB), 
	  .DDRA		                  (DDR_Addr),
	  .DDRBA		                (DDR_BankAddr),
	  .DDRCASB		              (DDR_CAS_n),
	  .DDRCKE		                (DDR_CKE),
	  .DDRCKN		                (DDR_Clk_n),
	  .DDRCKP		                (DDR_Clk),
	  .DDRCSB		                (DDR_CS_n),
	  .DDRDM		                (DDR_DM),
	  .DDRDQ		                (DDR_DQ),
	  .DDRDQSN		              (DDR_DQS_n),
	  .DDRDQSP		              (DDR_DQS),
	  .DDRDRSTB                 (DDR_DRSTB),
	  .DDRODT		                (DDR_ODT),  
	  .DDRRASB		              (DDR_RAS_n),
	  .DDRVRN                   (DDR_VRN),
	  .DDRVRP                   (DDR_VRP),
	  .DDRWEB                   (DDR_WEB),

    // 2 x PS Master PL Slave General Purpose Axi3 ports
	  .MAXIGP0ARESETN	          (M_AXI_GP0_ARESET_n),
	  .MAXIGP0ARADDR	          (M_AXI_GP0_ARADDR),
	  .MAXIGP0ARBURST	          (M_AXI_GP0_ARBURST),
    .MAXIGP0ARCACHE	          (M_AXI_GP0_ARCACHE),
	  .MAXIGP0ARID	            (M_AXI_GP0_ARID),
	  .MAXIGP0ARLEN	            (M_AXI_GP0_ARLEN),
	  .MAXIGP0ARLOCK	          (M_AXI_GP0_ARLOCK),
	  .MAXIGP0ARPROT	          (M_AXI_GP0_ARPROT),
	  .MAXIGP0ARQOS	            (M_AXI_GP0_ARQOS),
	  .MAXIGP0ARSIZE	          (M_AXI_GP0_ARSIZE),
	  .MAXIGP0ARVALID	          (M_AXI_GP0_ARVALID),
	  .MAXIGP0AWADDR	          (M_AXI_GP0_AWADDR),
	  .MAXIGP0AWBURST	          (M_AXI_GP0_AWBURST),
	  .MAXIGP0AWCACHE	          (M_AXI_GP0_AWCACHE),
	  .MAXIGP0AWID	            (M_AXI_GP0_AWID),
	  .MAXIGP0AWLEN	            (M_AXI_GP0_AWLEN),
	  .MAXIGP0AWLOCK	          (M_AXI_GP0_AWLOCK),
	  .MAXIGP0AWPROT	          (M_AXI_GP0_AWPROT),
	  .MAXIGP0AWQOS	            (M_AXI_GP0_AWQOS),
	  .MAXIGP0AWSIZE	          (M_AXI_GP0_AWSIZE),
	  .MAXIGP0AWVALID	          (M_AXI_GP0_AWVALID),
	  .MAXIGP0BREADY	          (M_AXI_GP0_BREADY),
	  .MAXIGP0RREADY	          (M_AXI_GP0_RREADY),
	  .MAXIGP0WDATA	            (M_AXI_GP0_WDATA),
	  .MAXIGP0WID	              (M_AXI_GP0_WID),
	  .MAXIGP0WLAST	            (M_AXI_GP0_WLAST),
	  .MAXIGP0WSTRB	            (M_AXI_GP0_WSTRB),
	  .MAXIGP0WVALID	          (M_AXI_GP0_WVALID),
	  .MAXIGP0ACLK	            (M_AXI_GP0_ACLK),
	  .MAXIGP0ARREADY	          (M_AXI_GP0_ARREADY),
	  .MAXIGP0AWREADY	          (M_AXI_GP0_AWREADY),
	  .MAXIGP0BID	              (M_AXI_GP0_BID),
	  .MAXIGP0BRESP	            (M_AXI_GP0_BRESP),
	  .MAXIGP0BVALID	          (M_AXI_GP0_BVALID),
	  .MAXIGP0RDATA	            (M_AXI_GP0_RDATA),
	  .MAXIGP0RID	              (M_AXI_GP0_RID),
	  .MAXIGP0RLAST	            (M_AXI_GP0_RLAST),
	  .MAXIGP0RRESP	            (M_AXI_GP0_RRESP),
	  .MAXIGP0RVALID	          (M_AXI_GP0_RVALID),
	  .MAXIGP0WREADY	          (M_AXI_GP0_WREADY),

	  .MAXIGP1ARESETN	          (M_AXI_GP1_ARESET_n),
	  .MAXIGP1ARADDR	          (M_AXI_GP1_ARADDR),
	  .MAXIGP1ARBURST	          (M_AXI_GP1_ARBURST),
	  .MAXIGP1ARCACHE	          (M_AXI_GP1_ARCACHE),
	  .MAXIGP1ARID	            (M_AXI_GP1_ARID),
	  .MAXIGP1ARLEN	            (M_AXI_GP1_ARLEN),
	  .MAXIGP1ARLOCK	          (M_AXI_GP1_ARLOCK),
	  .MAXIGP1ARPROT	          (M_AXI_GP1_ARPROT),
	  .MAXIGP1ARQOS	            (M_AXI_GP1_ARQOS),
	  .MAXIGP1ARSIZE	          (M_AXI_GP1_ARSIZE),
	  .MAXIGP1ARVALID	          (M_AXI_GP1_ARVALID),
	  .MAXIGP1AWADDR	          (M_AXI_GP1_AWADDR),
	  .MAXIGP1AWBURST	          (M_AXI_GP1_AWBURST),
	  .MAXIGP1AWCACHE	          (M_AXI_GP1_AWCACHE),
	  .MAXIGP1AWID	            (M_AXI_GP1_AWID),
	  .MAXIGP1AWLEN	            (M_AXI_GP1_AWLEN),
	  .MAXIGP1AWLOCK	          (M_AXI_GP1_AWLOCK),
	  .MAXIGP1AWPROT	          (M_AXI_GP1_AWPROT),
	  .MAXIGP1AWQOS	            (M_AXI_GP1_AWQOS),
	  .MAXIGP1AWSIZE	          (M_AXI_GP1_AWSIZE),
	  .MAXIGP1AWVALID	          (M_AXI_GP1_AWVALID),
	  .MAXIGP1BREADY	          (M_AXI_GP1_BREADY),
	  .MAXIGP1RREADY	          (M_AXI_GP1_RREADY),
	  .MAXIGP1WDATA	            (M_AXI_GP1_WDATA),
	  .MAXIGP1WID	              (M_AXI_GP1_WID),
	  .MAXIGP1WLAST	            (M_AXI_GP1_WLAST),
	  .MAXIGP1WSTRB	            (M_AXI_GP1_WSTRB),
	  .MAXIGP1WVALID	          (M_AXI_GP1_WVALID),
	  .MAXIGP1ACLK	            (M_AXI_GP1_ACLK),
	  .MAXIGP1ARREADY	          (M_AXI_GP1_ARREADY),
	  .MAXIGP1AWREADY	          (M_AXI_GP1_AWREADY),
	  .MAXIGP1BID	              (M_AXI_GP1_BID),
	  .MAXIGP1BRESP	            (M_AXI_GP1_BRESP),
	  .MAXIGP1BVALID	          (M_AXI_GP1_BVALID),
	  .MAXIGP1RDATA	            (M_AXI_GP1_RDATA),
	  .MAXIGP1RID	              (M_AXI_GP1_RID),
	  .MAXIGP1RLAST	            (M_AXI_GP1_RLAST),
	  .MAXIGP1RRESP	            (M_AXI_GP1_RRESP),
	  .MAXIGP1RVALID	          (M_AXI_GP1_RVALID),
	  .MAXIGP1WREADY	          (M_AXI_GP1_WREADY),  

    // 2 x PS Slave PL Master General Purpose Axi3 ports
	  .SAXIGP0ARESETN	          (S_AXI_GP0_ARESET_n),
	  .SAXIGP0ARREADY	          (S_AXI_GP0_ARREADY),
	  .SAXIGP0AWREADY	          (S_AXI_GP0_AWREADY),
	  .SAXIGP0BID	              (S_AXI_GP0_BID),
	  .SAXIGP0BRESP	            (S_AXI_GP0_BRESP),
	  .SAXIGP0BVALID	          (S_AXI_GP0_BVALID),
	  .SAXIGP0RDATA	            (S_AXI_GP0_RDATA),
	  .SAXIGP0RID	              (S_AXI_GP0_RID),
	  .SAXIGP0RLAST	            (S_AXI_GP0_RLAST),
	  .SAXIGP0RRESP	            (S_AXI_GP0_RRESP),
	  .SAXIGP0RVALID	          (S_AXI_GP0_RVALID),
	  .SAXIGP0WREADY	          (S_AXI_GP0_WREADY),
	  .SAXIGP0ACLK              (S_AXI_GP0_ACLK),
	  .SAXIGP0ARADDR            (S_AXI_GP0_ARADDR),
	  .SAXIGP0ARBURST           (S_AXI_GP0_ARBURST),
	  .SAXIGP0ARCACHE           (S_AXI_GP0_ARCACHE),
	  .SAXIGP0ARID              (S_AXI_GP0_ARID),
	  .SAXIGP0ARLEN             (S_AXI_GP0_ARLEN),
	  .SAXIGP0ARLOCK            (S_AXI_GP0_ARLOCK),
	  .SAXIGP0ARPROT            (S_AXI_GP0_ARPROT),
	  .SAXIGP0ARQOS             (S_AXI_GP0_ARQOS),
	  .SAXIGP0ARSIZE            (S_AXI_GP0_ARSIZE),
	  .SAXIGP0ARVALID           (S_AXI_GP0_ARVALID),
	  .SAXIGP0AWADDR            (S_AXI_GP0_AWADDR),
	  .SAXIGP0AWBURST           (S_AXI_GP0_AWBURST),
	  .SAXIGP0AWCACHE           (S_AXI_GP0_AWCACHE),
	  .SAXIGP0AWID              (S_AXI_GP0_AWID),
	  .SAXIGP0AWLEN             (S_AXI_GP0_AWLEN),
	  .SAXIGP0AWLOCK            (S_AXI_GP0_AWLOCK),
	  .SAXIGP0AWPROT            (S_AXI_GP0_AWPROT),
	  .SAXIGP0AWQOS             (S_AXI_GP0_AWQOS),
	  .SAXIGP0AWSIZE            (S_AXI_GP0_AWSIZE),
	  .SAXIGP0AWVALID           (S_AXI_GP0_AWVALID),
	  .SAXIGP0BREADY            (S_AXI_GP0_BREADY),
	  .SAXIGP0RREADY            (S_AXI_GP0_RREADY),
	  .SAXIGP0WDATA             (S_AXI_GP0_WDATA),
	  .SAXIGP0WID               (S_AXI_GP0_WID),
	  .SAXIGP0WLAST             (S_AXI_GP0_WLAST),
	  .SAXIGP0WSTRB             (S_AXI_GP0_WSTRB),
	  .SAXIGP0WVALID            (S_AXI_GP0_WVALID),

	  .SAXIGP1ARESETN	          (S_AXI_GP1_ARESET_n),
	  .SAXIGP1ARREADY	          (S_AXI_GP1_ARREADY),
	  .SAXIGP1AWREADY	          (S_AXI_GP1_AWREADY),
	  .SAXIGP1BID	              (S_AXI_GP1_BID),
	  .SAXIGP1BRESP	            (S_AXI_GP1_BRESP),
	  .SAXIGP1BVALID	          (S_AXI_GP1_BVALID),
	  .SAXIGP1RDATA	            (S_AXI_GP1_RDATA),
	  .SAXIGP1RID	              (S_AXI_GP1_RID),
	  .SAXIGP1RLAST	            (S_AXI_GP1_RLAST),
	  .SAXIGP1RRESP	            (S_AXI_GP1_RRESP),
	  .SAXIGP1RVALID	          (S_AXI_GP1_RVALID),
	  .SAXIGP1WREADY	          (S_AXI_GP1_WREADY),
	  .SAXIGP1ACLK	            (S_AXI_GP1_ACLK),
	  .SAXIGP1ARADDR	          (S_AXI_GP1_ARADDR),
	  .SAXIGP1ARBURST	          (S_AXI_GP1_ARBURST),
	  .SAXIGP1ARCACHE	          (S_AXI_GP1_ARCACHE),
	  .SAXIGP1ARID	            (S_AXI_GP1_ARID),
	  .SAXIGP1ARLEN	            (S_AXI_GP1_ARLEN),
	  .SAXIGP1ARLOCK	          (S_AXI_GP1_ARLOCK),
	  .SAXIGP1ARPROT	          (S_AXI_GP1_ARPROT),
	  .SAXIGP1ARQOS	            (S_AXI_GP1_ARQOS),
	  .SAXIGP1ARSIZE	          (S_AXI_GP1_ARSIZE),
	  .SAXIGP1ARVALID	          (S_AXI_GP1_ARVALID),
	  .SAXIGP1AWADDR	          (S_AXI_GP1_AWADDR),
	  .SAXIGP1AWBURST	          (S_AXI_GP1_AWBURST),
	  .SAXIGP1AWCACHE	          (S_AXI_GP1_AWCACHE),
	  .SAXIGP1AWID	            (S_AXI_GP1_AWID),
	  .SAXIGP1AWLEN	            (S_AXI_GP1_AWLEN),
	  .SAXIGP1AWLOCK	          (S_AXI_GP1_AWLOCK),
	  .SAXIGP1AWPROT	          (S_AXI_GP1_AWPROT),
	  .SAXIGP1AWQOS	            (S_AXI_GP1_AWQOS),
	  .SAXIGP1AWSIZE	          (S_AXI_GP1_AWSIZE),
	  .SAXIGP1AWVALID	          (S_AXI_GP1_AWVALID),
	  .SAXIGP1BREADY	          (S_AXI_GP1_BREADY),
	  .SAXIGP1RREADY	          (S_AXI_GP1_RREADY),
	  .SAXIGP1WDATA	            (S_AXI_GP1_WDATA),
	  .SAXIGP1WID	              (S_AXI_GP1_WID),
	  .SAXIGP1WLAST	            (S_AXI_GP1_WLAST),
	  .SAXIGP1WSTRB	            (S_AXI_GP1_WSTRB),
	  .SAXIGP1WVALID	          (S_AXI_GP1_WVALID),  

    // 1x PS Slave PL Master ACP Axi3 port
	  .SAXIACPARESETN	          (S_AXI_ACP_ARESET_n),
	  .SAXIACPARREADY	          (S_AXI_ACP_ARREADY),
	  .SAXIACPAWREADY	          (S_AXI_ACP_AWREADY),
	  .SAXIACPBID	              (S_AXI_ACP_BID),
	  .SAXIACPBRESP	            (S_AXI_ACP_BRESP),
	  .SAXIACPBVALID	          (S_AXI_ACP_BVALID),
	  .SAXIACPRDATA	            (S_AXI_ACP_RDATA),
	  .SAXIACPRID	              (S_AXI_ACP_RID),
	  .SAXIACPRLAST	            (S_AXI_ACP_RLAST),
	  .SAXIACPRRESP	            (S_AXI_ACP_RRESP),
	  .SAXIACPRVALID	          (S_AXI_ACP_RVALID),
	  .SAXIACPWREADY	          (S_AXI_ACP_WREADY),
	  .SAXIACPACLK	            (S_AXI_ACP_ACLK),
	  .SAXIACPARADDR	          (S_AXI_ACP_ARADDR),
	  .SAXIACPARBURST	          (S_AXI_ACP_ARBURST),
	  .SAXIACPARCACHE	          (S_AXI_ACP_ARCACHE),
	  .SAXIACPARID	            (S_AXI_ACP_ARID),
	  .SAXIACPARLEN	            (S_AXI_ACP_ARLEN),
	  .SAXIACPARLOCK	          (S_AXI_ACP_ARLOCK),
	  .SAXIACPARPROT	          (S_AXI_ACP_ARPROT),
	  .SAXIACPARQOS	            (S_AXI_ACP_ARQOS),
	  .SAXIACPARSIZE	          (S_AXI_ACP_ARSIZE),
	  .SAXIACPARVALID	          (S_AXI_ACP_ARVALID),
	  .SAXIACPAWADDR	          (S_AXI_ACP_AWADDR),
	  .SAXIACPAWBURST	          (S_AXI_ACP_AWBURST),
	  .SAXIACPAWCACHE	          (S_AXI_ACP_AWCACHE),
	  .SAXIACPAWID	            (S_AXI_ACP_AWID),
	  .SAXIACPAWLEN	            (S_AXI_ACP_AWLEN),
	  .SAXIACPAWLOCK	          (S_AXI_ACP_AWLOCK),
	  .SAXIACPAWPROT	          (S_AXI_ACP_AWPROT),
	  .SAXIACPAWQOS	            (S_AXI_ACP_AWQOS),
	  .SAXIACPAWSIZE	          (S_AXI_ACP_AWSIZE),
	  .SAXIACPAWVALID	          (S_AXI_ACP_AWVALID),
	  .SAXIACPBREADY	          (S_AXI_ACP_BREADY),
	  .SAXIACPRREADY	          (S_AXI_ACP_RREADY),
	  .SAXIACPWDATA	            (S_AXI_ACP_WDATA),
	  .SAXIACPWID	              (S_AXI_ACP_WID),
	  .SAXIACPWLAST	            (S_AXI_ACP_WLAST),
	  .SAXIACPWSTRB	            (S_AXI_ACP_WSTRB),
	  .SAXIACPWVALID	          (S_AXI_ACP_WVALID),
    .SAXIACPARUSER            (S_AXI_ACP_ARUSER),
    .SAXIACPAWUSER            (S_AXI_ACP_AWUSER),

    // 4x PS Slave PL Master High Performance Axi3 port
	  .SAXIHP0ARESETN	          (S_AXI_HP0_ARESETN),
	  .SAXIHP0ARREADY	          (S_AXI_HP0_ARREADY),
	  .SAXIHP0AWREADY	          (S_AXI_HP0_AWREADY),
	  .SAXIHP0BID	              (S_AXI_HP0_BID),
	  .SAXIHP0BRESP	            (S_AXI_HP0_BRESP),
	  .SAXIHP0BVALID	          (S_AXI_HP0_BVALID),
	  .SAXIHP0RACOUNT           (S_AXI_HP0_RACOUNT),
	  .SAXIHP0RCOUNT	          (S_AXI_HP0_RCOUNT),
	  .SAXIHP0RDATA	            (S_AXI_HP0_RDATA),
	  .SAXIHP0RID	              (S_AXI_HP0_RID),
	  .SAXIHP0RLAST	            (S_AXI_HP0_RLAST),
	  .SAXIHP0RRESP	            (S_AXI_HP0_RRESP),
	  .SAXIHP0RVALID	          (S_AXI_HP0_RVALID),
	  .SAXIHP0WCOUNT	          (S_AXI_HP0_WCOUNT),
	  .SAXIHP0WACOUNT           (S_AXI_HP0_WACOUNT),  
	  .SAXIHP0WREADY	          (S_AXI_HP0_WREADY),
	  .SAXIHP0ACLK              (S_AXI_HP0_ACLK),
	  .SAXIHP0ARADDR            (S_AXI_HP0_ARADDR),
	  .SAXIHP0ARBURST           (S_AXI_HP0_ARBURST),
	  .SAXIHP0ARCACHE           (S_AXI_HP0_ARCACHE),
	  .SAXIHP0ARID              (S_AXI_HP0_ARID),
	  .SAXIHP0ARLEN             (S_AXI_HP0_ARLEN),
	  .SAXIHP0ARLOCK            (S_AXI_HP0_ARLOCK),
	  .SAXIHP0ARPROT            (S_AXI_HP0_ARPROT),
	  .SAXIHP0ARQOS             (S_AXI_HP0_ARQOS),
	  .SAXIHP0ARSIZE            (S_AXI_HP0_ARSIZE),
	  .SAXIHP0ARVALID           (S_AXI_HP0_ARVALID),
	  .SAXIHP0AWADDR            (S_AXI_HP0_AWADDR),
	  .SAXIHP0AWBURST           (S_AXI_HP0_AWBURST),
	  .SAXIHP0AWCACHE           (S_AXI_HP0_AWCACHE),
	  .SAXIHP0AWID              (S_AXI_HP0_AWID),
	  .SAXIHP0AWLEN             (S_AXI_HP0_AWLEN),
	  .SAXIHP0AWLOCK            (S_AXI_HP0_AWLOCK),
	  .SAXIHP0AWPROT            (S_AXI_HP0_AWPROT),
	  .SAXIHP0AWQOS             (S_AXI_HP0_AWQOS),
	  .SAXIHP0AWSIZE            (S_AXI_HP0_AWSIZE),
	  .SAXIHP0AWVALID           (S_AXI_HP0_AWVALID),
	  .SAXIHP0BREADY            (S_AXI_HP0_BREADY),
	  .SAXIHP0RDISSUECAP1EN     (S_AXI_HP0_RDISSUECAP1_EN),
	  .SAXIHP0RREADY            (S_AXI_HP0_RREADY),
	  .SAXIHP0WDATA             (S_AXI_HP0_WDATA),
	  .SAXIHP0WID               (S_AXI_HP0_WID),
	  .SAXIHP0WLAST             (S_AXI_HP0_WLAST),
	  .SAXIHP0WRISSUECAP1EN     (S_AXI_HP0_WRISSUECAP1_EN),
	  .SAXIHP0WSTRB             (S_AXI_HP0_WSTRB),
	  .SAXIHP0WVALID            (S_AXI_HP0_WVALID),


	  .SAXIHP1ACLK              (S_AXI_HP1_ACLK),
	  .SAXIHP1ARADDR            (S_AXI_HP1_ARADDR),
	  .SAXIHP1ARBURST           (S_AXI_HP1_ARBURST),
	  .SAXIHP1ARCACHE           (S_AXI_HP1_ARCACHE),
	  .SAXIHP1ARID              (S_AXI_HP1_ARID),
	  .SAXIHP1ARLEN             (S_AXI_HP1_ARLEN),
	  .SAXIHP1ARLOCK            (S_AXI_HP1_ARLOCK),
	  .SAXIHP1ARPROT            (S_AXI_HP1_ARPROT),
	  .SAXIHP1ARQOS             (S_AXI_HP1_ARQOS),
	  .SAXIHP1ARSIZE            (S_AXI_HP1_ARSIZE),
	  .SAXIHP1ARVALID           (S_AXI_HP1_ARVALID),
	  .SAXIHP1AWADDR            (S_AXI_HP1_AWADDR),
	  .SAXIHP1AWBURST           (S_AXI_HP1_AWBURST),
	  .SAXIHP1AWCACHE           (S_AXI_HP1_AWCACHE),
	  .SAXIHP1AWID              (S_AXI_HP1_AWID),
	  .SAXIHP1AWLEN             (S_AXI_HP1_AWLEN),
	  .SAXIHP1AWLOCK            (S_AXI_HP1_AWLOCK),
	  .SAXIHP1AWPROT            (S_AXI_HP1_AWPROT),
	  .SAXIHP1AWQOS             (S_AXI_HP1_AWQOS),
	  .SAXIHP1AWSIZE            (S_AXI_HP1_AWSIZE),
	  .SAXIHP1AWVALID           (S_AXI_HP1_AWVALID),
	  .SAXIHP1BREADY            (S_AXI_HP1_BREADY),
	  .SAXIHP1RDISSUECAP1EN     (S_AXI_HP1_RDISSUECAP1_EN),
	  .SAXIHP1RREADY            (S_AXI_HP1_RREADY),
	  .SAXIHP1WDATA             (S_AXI_HP1_WDATA),
	  .SAXIHP1WID               (S_AXI_HP1_WID),
	  .SAXIHP1WLAST             (S_AXI_HP1_WLAST),
	  .SAXIHP1WRISSUECAP1EN     (S_AXI_HP1_WRISSUECAP1_EN),
	  .SAXIHP1WSTRB             (S_AXI_HP1_WSTRB),
	  .SAXIHP1WVALID            (S_AXI_HP1_WVALID),
	  .SAXIHP1ARESETN	          (S_AXI_HP1_ARESETN),
	  .SAXIHP1ARREADY	          (S_AXI_HP1_ARREADY),
	  .SAXIHP1AWREADY	          (S_AXI_HP1_AWREADY),
	  .SAXIHP1BID	              (S_AXI_HP1_BID),
	  .SAXIHP1BRESP	            (S_AXI_HP1_BRESP),
	  .SAXIHP1BVALID	          (S_AXI_HP1_BVALID),
	  .SAXIHP1RACOUNT	          (S_AXI_HP1_RACOUNT),  
	  .SAXIHP1RCOUNT	          (S_AXI_HP1_RCOUNT),
	  .SAXIHP1RDATA	            (S_AXI_HP1_RDATA),
	  .SAXIHP1RID	              (S_AXI_HP1_RID),
	  .SAXIHP1RLAST	            (S_AXI_HP1_RLAST),
	  .SAXIHP1RRESP	            (S_AXI_HP1_RRESP),
	  .SAXIHP1RVALID	          (S_AXI_HP1_RVALID),
	  .SAXIHP1WACOUNT	          (S_AXI_HP1_WACOUNT),  
	  .SAXIHP1WCOUNT	          (S_AXI_HP1_WCOUNT),
	  .SAXIHP1WREADY	          (S_AXI_HP1_WREADY),

	  .SAXIHP2ARESETN	          (S_AXI_HP2_ARESET_n),
	  .SAXIHP2ARREADY	          (S_AXI_HP2_ARREADY),
	  .SAXIHP2AWREADY	          (S_AXI_HP2_AWREADY),
	  .SAXIHP2BID	              (S_AXI_HP2_BID),
	  .SAXIHP2BRESP	            (S_AXI_HP2_BRESP),
	  .SAXIHP2BVALID	          (S_AXI_HP2_BVALID),
	  .SAXIHP2RACOUNT	          (S_AXI_HP2_RACOUNT),  
	  .SAXIHP2RCOUNT	          (S_AXI_HP2_RCOUNT),
	  .SAXIHP2RDATA	            (S_AXI_HP2_RDATA),
	  .SAXIHP2RID	              (S_AXI_HP2_RID),
	  .SAXIHP2RLAST	            (S_AXI_HP2_RLAST),
	  .SAXIHP2RRESP	            (S_AXI_HP2_RRESP),
	  .SAXIHP2RVALID	          (S_AXI_HP2_RVALID),
	  .SAXIHP2WACOUNT	          (S_AXI_HP2_WACOUNT),  
	  .SAXIHP2WCOUNT	          (S_AXI_HP2_WCOUNT),
	  .SAXIHP2WREADY	          (S_AXI_HP2_WREADY),
	  .SAXIHP2ACLK              (S_AXI_HP2_ACLK),
	  .SAXIHP2ARADDR            (S_AXI_HP2_ARADDR),
	  .SAXIHP2ARBURST           (S_AXI_HP2_ARBURST),
	  .SAXIHP2ARCACHE           (S_AXI_HP2_ARCACHE),
	  .SAXIHP2ARID              (S_AXI_HP2_ARID),
	  .SAXIHP2ARLEN             (S_AXI_HP2_ARLEN),
	  .SAXIHP2ARLOCK            (S_AXI_HP2_ARLOCK),
	  .SAXIHP2ARPROT            (S_AXI_HP2_ARPROT),
	  .SAXIHP2ARQOS             (S_AXI_HP2_ARQOS),
	  .SAXIHP2ARSIZE            (S_AXI_HP2_ARSIZE),
	  .SAXIHP2ARVALID           (S_AXI_HP2_ARVALID),
	  .SAXIHP2AWADDR            (S_AXI_HP2_AWADDR),
	  .SAXIHP2AWBURST           (S_AXI_HP2_AWBURST),
	  .SAXIHP2AWCACHE           (S_AXI_HP2_AWCACHE),
	  .SAXIHP2AWID              (S_AXI_HP2_AWID),
	  .SAXIHP2AWLEN             (S_AXI_HP2_AWLEN),
	  .SAXIHP2AWLOCK            (S_AXI_HP2_AWLOCK),
	  .SAXIHP2AWPROT            (S_AXI_HP2_AWPROT),
	  .SAXIHP2AWQOS             (S_AXI_HP2_AWQOS),
	  .SAXIHP2AWSIZE            (S_AXI_HP2_AWSIZE),
	  .SAXIHP2AWVALID           (S_AXI_HP2_AWVALID),
	  .SAXIHP2BREADY            (S_AXI_HP2_BREADY),
	  .SAXIHP2RDISSUECAP1EN     (S_AXI_HP2_RDISSUECAP1_EN),
	  .SAXIHP2RREADY            (S_AXI_HP2_RREADY),
	  .SAXIHP2WDATA             (S_AXI_HP2_WDATA),
	  .SAXIHP2WID               (S_AXI_HP2_WID),
	  .SAXIHP2WLAST             (S_AXI_HP2_WLAST),
	  .SAXIHP2WRISSUECAP1EN     (S_AXI_HP2_WRISSUECAP1_EN),
	  .SAXIHP2WSTRB             (S_AXI_HP2_WSTRB),
	  .SAXIHP2WVALID            (S_AXI_HP2_WVALID),  

	  .SAXIHP3ARESETN	          (S_AXI_HP3_ARESET_n),
	  .SAXIHP3ARREADY	          (S_AXI_HP3_ARREADY),
	  .SAXIHP3AWREADY	          (S_AXI_HP3_AWREADY),
	  .SAXIHP3BID	              (S_AXI_HP3_BID),
	  .SAXIHP3BRESP	            (S_AXI_HP3_BRESP),
	  .SAXIHP3BVALID	          (S_AXI_HP3_BVALID),
	  .SAXIHP3RACOUNT	          (S_AXI_HP3_RACOUNT),    
	  .SAXIHP3RCOUNT	          (S_AXI_HP3_RCOUNT),
	  .SAXIHP3RDATA	            (S_AXI_HP3_RDATA),
	  .SAXIHP3RID	              (S_AXI_HP3_RID),
	  .SAXIHP3RLAST	            (S_AXI_HP3_RLAST),
	  .SAXIHP3RRESP	            (S_AXI_HP3_RRESP),
	  .SAXIHP3RVALID	          (S_AXI_HP3_RVALID),
	  .SAXIHP3WCOUNT	          (S_AXI_HP3_WCOUNT),
	  .SAXIHP3WACOUNT	          (S_AXI_HP3_WACOUNT),    
	  .SAXIHP3WREADY	          (S_AXI_HP3_WREADY), 
	  .SAXIHP3ACLK              (S_AXI_HP3_ACLK),
	  .SAXIHP3ARADDR            (S_AXI_HP3_ARADDR),
	  .SAXIHP3ARBURST           (S_AXI_HP3_ARBURST),
	  .SAXIHP3ARCACHE           (S_AXI_HP3_ARCACHE),
	  .SAXIHP3ARID              (S_AXI_HP3_ARID),
	  .SAXIHP3ARLEN             (S_AXI_HP3_ARLEN),
	  .SAXIHP3ARLOCK            (S_AXI_HP3_ARLOCK),
	  .SAXIHP3ARPROT            (S_AXI_HP3_ARPROT),
	  .SAXIHP3ARQOS             (S_AXI_HP3_ARQOS),
	  .SAXIHP3ARSIZE            (S_AXI_HP3_ARSIZE),
	  .SAXIHP3ARVALID           (S_AXI_HP3_ARVALID),
	  .SAXIHP3AWADDR            (S_AXI_HP3_AWADDR),
	  .SAXIHP3AWBURST           (S_AXI_HP3_AWBURST),
	  .SAXIHP3AWCACHE           (S_AXI_HP3_AWCACHE),
	  .SAXIHP3AWID              (S_AXI_HP3_AWID),
	  .SAXIHP3AWLEN             (S_AXI_HP3_AWLEN),
	  .SAXIHP3AWLOCK            (S_AXI_HP3_AWLOCK),
	  .SAXIHP3AWPROT            (S_AXI_HP3_AWPROT),
	  .SAXIHP3AWQOS             (S_AXI_HP3_AWQOS),
	  .SAXIHP3AWSIZE            (S_AXI_HP3_AWSIZE),
	  .SAXIHP3AWVALID           (S_AXI_HP3_AWVALID),
	  .SAXIHP3BREADY            (S_AXI_HP3_BREADY),
	  .SAXIHP3RDISSUECAP1EN     (S_AXI_HP3_RDISSUECAP1_EN),
	  .SAXIHP3RREADY            (S_AXI_HP3_RREADY),
	  .SAXIHP3WDATA             (S_AXI_HP3_WDATA),
	  .SAXIHP3WID               (S_AXI_HP3_WID),
	  .SAXIHP3WLAST             (S_AXI_HP3_WLAST),
	  .SAXIHP3WRISSUECAP1EN     (S_AXI_HP3_WRISSUECAP1_EN),
	  .SAXIHP3WSTRB             (S_AXI_HP3_WSTRB),
	  .SAXIHP3WVALID            (S_AXI_HP3_WVALID) 
	);

endmodule
